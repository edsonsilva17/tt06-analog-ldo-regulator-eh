magic
tech sky130A
timestamp 1712983369
<< metal1 >>
rect -115 13310 0 13410
rect 4550 9770 4565 9870
rect 7600 9770 7715 9870
rect -115 8090 0 8190
rect 1250 8180 4775 8190
rect 1250 8100 4685 8180
rect 4765 8100 4775 8180
rect 1250 8090 4775 8100
rect 7585 6105 7700 6205
rect 4575 4570 4655 4645
rect 7600 4570 7700 4580
rect 4575 4490 7700 4570
rect 7600 4480 7700 4490
<< via1 >>
rect 4685 8100 4765 8180
<< metal2 >>
rect 4675 8180 7465 8190
rect 4675 8100 4685 8180
rect 4765 8100 7465 8180
rect 4675 8090 7465 8100
use cell  x1
timestamp 1712944235
transform 1 0 450 0 1 8000
box -450 -7700 4100 5410
use LDO  x2
timestamp 1712939325
transform 1 0 4565 0 1 4395
box 0 250 3035 5475
<< labels >>
flabel metal1 -115 13310 -15 13410 0 FreeSans 128 0 0 0 top_in
port 0 nsew
flabel metal1 -115 8090 -15 8190 0 FreeSans 128 0 0 0 top_gnd
port 1 nsew
flabel metal1 7615 9770 7715 9870 0 FreeSans 128 0 0 0 top_out
port 4 nsew
flabel metal1 7600 6105 7700 6205 0 FreeSans 128 0 0 0 top_ref
port 3 nsew
flabel metal1 7600 4480 7700 4580 0 FreeSans 128 0 0 0 top_ibias
port 2 nsew
<< end >>
