magic
tech sky130A
magscale 1 2
timestamp 1712843110
<< metal3 >>
rect -3150 9372 3149 9400
rect -3150 3228 3065 9372
rect 3129 3228 3149 9372
rect -3150 3200 3149 3228
rect -3150 3072 3149 3100
rect -3150 -3072 3065 3072
rect 3129 -3072 3149 3072
rect -3150 -3100 3149 -3072
rect -3150 -3228 3149 -3200
rect -3150 -9372 3065 -3228
rect 3129 -9372 3149 -3228
rect -3150 -9400 3149 -9372
<< via3 >>
rect 3065 3228 3129 9372
rect 3065 -3072 3129 3072
rect 3065 -9372 3129 -3228
<< mimcap >>
rect -3050 9260 2950 9300
rect -3050 3340 -3010 9260
rect 2910 3340 2950 9260
rect -3050 3300 2950 3340
rect -3050 2960 2950 3000
rect -3050 -2960 -3010 2960
rect 2910 -2960 2950 2960
rect -3050 -3000 2950 -2960
rect -3050 -3340 2950 -3300
rect -3050 -9260 -3010 -3340
rect 2910 -9260 2950 -3340
rect -3050 -9300 2950 -9260
<< mimcapcontact >>
rect -3010 3340 2910 9260
rect -3010 -2960 2910 2960
rect -3010 -9260 2910 -3340
<< metal4 >>
rect -102 9261 2 9450
rect 3018 9388 3122 9450
rect 3018 9372 3145 9388
rect -3011 9260 2911 9261
rect -3011 3340 -3010 9260
rect 2910 3340 2911 9260
rect -3011 3339 2911 3340
rect -102 2961 2 3339
rect 3018 3228 3065 9372
rect 3129 3228 3145 9372
rect 3018 3212 3145 3228
rect 3018 3088 3122 3212
rect 3018 3072 3145 3088
rect -3011 2960 2911 2961
rect -3011 -2960 -3010 2960
rect 2910 -2960 2911 2960
rect -3011 -2961 2911 -2960
rect -102 -3339 2 -2961
rect 3018 -3072 3065 3072
rect 3129 -3072 3145 3072
rect 3018 -3088 3145 -3072
rect 3018 -3212 3122 -3088
rect 3018 -3228 3145 -3212
rect -3011 -3340 2911 -3339
rect -3011 -9260 -3010 -3340
rect 2910 -9260 2911 -3340
rect -3011 -9261 2911 -9260
rect -102 -9450 2 -9261
rect 3018 -9372 3065 -3228
rect 3129 -9372 3145 -3228
rect 3018 -9388 3145 -9372
rect 3018 -9450 3122 -9388
<< properties >>
string FIXED_BBOX -3150 3200 3050 9400
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.0 l 30.0 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
