magic
tech sky130A
magscale 1 2
timestamp 1712930611
<< metal1 >>
rect 5220 500 5420 530
rect -150 480 5420 500
rect -150 370 5060 480
rect 5160 370 5420 480
rect -150 350 5420 370
rect -150 -710 10 350
rect 5220 330 5420 350
rect 1580 170 5400 190
rect 1580 60 5260 170
rect 5380 60 5400 170
rect 1580 40 5400 60
rect 4160 -60 4170 -50
rect 1770 -130 4170 -60
rect 4160 -140 4170 -130
rect 4260 -140 4270 -50
rect -150 -860 3280 -710
rect 5220 -820 5420 -770
rect 4260 -920 5420 -820
rect -150 -1180 3540 -1030
rect 4260 -1180 4360 -920
rect 5220 -970 5420 -920
rect -150 -1310 40 -1180
rect -150 -2110 10 -1310
rect 190 -1360 3490 -1270
rect 1040 -1650 1130 -1360
rect 3980 -1500 4240 -1350
rect 4370 -1370 4890 -1350
rect 4370 -1480 4600 -1370
rect 4710 -1480 4890 -1370
rect 4370 -1500 4890 -1480
rect 5010 -1370 5400 -1350
rect 5010 -1480 5260 -1370
rect 5380 -1480 5400 -1370
rect 5010 -1500 5400 -1480
rect 1040 -1660 3490 -1650
rect 1040 -1730 1050 -1660
rect 1120 -1730 3490 -1660
rect 1040 -1740 3490 -1730
rect 3980 -1830 4060 -1500
rect 1430 -1980 4060 -1830
rect 4900 -1850 5000 -1660
rect 5240 -1780 5400 -1500
rect -170 -2140 30 -2110
rect -170 -2290 3274 -2140
rect 3980 -2270 4060 -1980
rect 4600 -1910 5000 -1850
rect 4600 -2270 4700 -1910
rect 4900 -2100 5000 -1910
rect 5220 -1980 5420 -1780
rect 5240 -2270 5400 -1980
rect -170 -2310 30 -2290
rect -150 -2960 10 -2310
rect 3980 -2420 4240 -2270
rect 4370 -2420 4890 -2270
rect 5010 -2420 5400 -2270
rect 4260 -2840 4360 -2580
rect 5220 -2840 5420 -2790
rect 4260 -2940 5420 -2840
rect -150 -3110 3534 -2960
rect 5220 -2990 5420 -2940
rect -170 -3270 30 -3240
rect -170 -3300 3280 -3270
rect -170 -3390 1040 -3300
rect 1130 -3390 3280 -3300
rect -170 -3420 3280 -3390
rect -170 -3440 30 -3420
rect 1040 -3510 1130 -3420
rect 1040 -3600 3490 -3510
<< via1 >>
rect 5060 370 5160 480
rect 5260 60 5380 170
rect 4170 -140 4260 -50
rect 4600 -1480 4710 -1370
rect 5260 -1480 5380 -1370
rect 1050 -1730 1120 -1660
rect 1040 -3390 1130 -3300
<< metal2 >>
rect 5060 480 5160 490
rect 5060 360 5160 370
rect 5240 170 5400 190
rect 5240 60 5260 170
rect 5380 60 5400 170
rect 4160 -50 4270 -40
rect 4160 -140 4170 -50
rect 4260 -140 4270 -50
rect 4160 -660 4270 -140
rect 4160 -770 4710 -660
rect 4600 -1370 4710 -770
rect 4600 -1490 4710 -1480
rect 5240 -1370 5400 60
rect 5240 -1480 5260 -1370
rect 5380 -1480 5400 -1370
rect 5240 -1500 5400 -1480
rect 1040 -1660 1130 -1650
rect 1040 -1730 1050 -1660
rect 1120 -1730 1130 -1660
rect 1040 -3300 1130 -1730
rect 1040 -3400 1130 -3390
<< via2 >>
rect 5060 370 5160 480
rect 4170 -140 4260 -50
<< metal3 >>
rect 5050 480 5170 485
rect 5050 370 5060 480
rect 5160 370 5170 480
rect 5050 365 5170 370
rect 4160 -50 4270 -45
rect 4160 -140 4170 -50
rect 4260 -140 4270 -50
rect 4160 -145 4270 -140
<< via3 >>
rect 5060 370 5160 480
rect 4170 -140 4260 -50
<< metal4 >>
rect 4160 -50 4270 1110
rect 5060 481 5160 890
rect 5059 480 5161 481
rect 5059 370 5060 480
rect 5160 370 5161 480
rect 5059 369 5161 370
rect 4160 -140 4170 -50
rect 4260 -140 4270 -50
rect 4160 -150 4270 -140
use sky130_fd_pr__cap_mim_m3_1_M5BWMD  XC1
timestamp 1712927986
transform 1 0 2710 0 1 3250
box -2450 -2400 2449 2400
use sky130_fd_pr__pfet_g5v0d10v5_4LQ75H  XM1
timestamp 1712930052
transform -1 0 4308 0 -1 -2343
box -308 -497 308 497
use sky130_fd_pr__pfet_g5v0d10v5_LMT75H  XM2
timestamp 1712930052
transform 1 0 4308 0 1 -1423
box -308 -497 308 497
use sky130_fd_pr__nfet_g5v0d10v5_RVNTYK  XM3
timestamp 1712930560
transform -1 0 4950 0 -1 -2830
box -278 -958 278 958
use sky130_fd_pr__nfet_g5v0d10v5_RMPAXK  XM4
timestamp 1712930560
transform 1 0 4950 0 1 -930
box -278 -958 278 958
use sky130_fd_pr__pfet_g5v0d10v5_FYUU4F  XM5
timestamp 1712928946
transform 1 0 2481 0 1 -2063
box -1261 -597 1261 597
use sky130_fd_pr__pfet_g5v0d10v5_C5553C  XM6
timestamp 1712928946
transform 1 0 1836 0 1 -943
box -1906 -597 1906 597
use sky130_fd_pr__nfet_g5v0d10v5_YCT7Q3  XM7
timestamp 1712930560
transform 1 0 2644 0 1 270
box -1102 -558 1102 558
use sky130_fd_pr__pfet_g5v0d10v5_FY4V4F  XM8
timestamp 1712930611
transform 1 0 2481 0 1 -3193
box -1261 -597 1261 597
<< labels >>
flabel metal1 -170 -2310 30 -2110 0 FreeSans 256 0 0 0 VDD
port 2 nsew
flabel metal1 -170 -3440 30 -3240 0 FreeSans 256 0 0 0 Ibias
port 4 nsew
flabel metal1 5220 -1980 5420 -1780 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 5220 330 5420 530 0 FreeSans 256 0 0 0 Vout
port 5 nsew
flabel metal1 5220 -970 5420 -770 0 FreeSans 256 0 0 0 Vip
port 1 nsew
flabel metal1 5220 -2990 5420 -2790 0 FreeSans 256 0 0 0 Vin
port 0 nsew
<< end >>
