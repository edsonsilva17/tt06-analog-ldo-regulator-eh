magic
tech sky130A
magscale 1 2
timestamp 1713034554
<< nwell >>
rect -1261 -597 1261 597
<< mvpmos >>
rect -1003 -300 -803 300
rect -745 -300 -545 300
rect -487 -300 -287 300
rect -229 -300 -29 300
rect 29 -300 229 300
rect 287 -300 487 300
rect 545 -300 745 300
rect 803 -300 1003 300
<< mvpdiff >>
rect -1061 288 -1003 300
rect -1061 -288 -1049 288
rect -1015 -288 -1003 288
rect -1061 -300 -1003 -288
rect -803 288 -745 300
rect -803 -288 -791 288
rect -757 -288 -745 288
rect -803 -300 -745 -288
rect -545 288 -487 300
rect -545 -288 -533 288
rect -499 -288 -487 288
rect -545 -300 -487 -288
rect -287 288 -229 300
rect -287 -288 -275 288
rect -241 -288 -229 288
rect -287 -300 -229 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 229 288 287 300
rect 229 -288 241 288
rect 275 -288 287 288
rect 229 -300 287 -288
rect 487 288 545 300
rect 487 -288 499 288
rect 533 -288 545 288
rect 487 -300 545 -288
rect 745 288 803 300
rect 745 -288 757 288
rect 791 -288 803 288
rect 745 -300 803 -288
rect 1003 288 1061 300
rect 1003 -288 1015 288
rect 1049 -288 1061 288
rect 1003 -300 1061 -288
<< mvpdiffc >>
rect -1049 -288 -1015 288
rect -791 -288 -757 288
rect -533 -288 -499 288
rect -275 -288 -241 288
rect -17 -288 17 288
rect 241 -288 275 288
rect 499 -288 533 288
rect 757 -288 791 288
rect 1015 -288 1049 288
<< mvnsubdiff >>
rect -1195 519 1195 531
rect -1195 485 -1087 519
rect 1087 485 1195 519
rect -1195 473 1195 485
rect -1195 423 -1137 473
rect -1195 -423 -1183 423
rect -1149 -423 -1137 423
rect 1137 423 1195 473
rect -1195 -473 -1137 -423
rect 1137 -423 1149 423
rect 1183 -423 1195 423
rect 1137 -473 1195 -423
rect -1195 -485 1195 -473
rect -1195 -519 -1087 -485
rect 1087 -519 1195 -485
rect -1195 -531 1195 -519
<< mvnsubdiffcont >>
rect -1087 485 1087 519
rect -1183 -423 -1149 423
rect 1149 -423 1183 423
rect -1087 -519 1087 -485
<< poly >>
rect -1003 381 -803 397
rect -1003 347 -987 381
rect -819 347 -803 381
rect -1003 300 -803 347
rect -745 381 -545 397
rect -745 347 -729 381
rect -561 347 -545 381
rect -745 300 -545 347
rect -487 381 -287 397
rect -487 347 -471 381
rect -303 347 -287 381
rect -487 300 -287 347
rect -229 381 -29 397
rect -229 347 -213 381
rect -45 347 -29 381
rect -229 300 -29 347
rect 29 381 229 397
rect 29 347 45 381
rect 213 347 229 381
rect 29 300 229 347
rect 287 381 487 397
rect 287 347 303 381
rect 471 347 487 381
rect 287 300 487 347
rect 545 381 745 397
rect 545 347 561 381
rect 729 347 745 381
rect 545 300 745 347
rect 803 381 1003 397
rect 803 347 819 381
rect 987 347 1003 381
rect 803 300 1003 347
rect -1003 -347 -803 -300
rect -1003 -381 -987 -347
rect -819 -381 -803 -347
rect -1003 -397 -803 -381
rect -745 -347 -545 -300
rect -745 -381 -729 -347
rect -561 -381 -545 -347
rect -745 -397 -545 -381
rect -487 -347 -287 -300
rect -487 -381 -471 -347
rect -303 -381 -287 -347
rect -487 -397 -287 -381
rect -229 -347 -29 -300
rect -229 -381 -213 -347
rect -45 -381 -29 -347
rect -229 -397 -29 -381
rect 29 -347 229 -300
rect 29 -381 45 -347
rect 213 -381 229 -347
rect 29 -397 229 -381
rect 287 -347 487 -300
rect 287 -381 303 -347
rect 471 -381 487 -347
rect 287 -397 487 -381
rect 545 -347 745 -300
rect 545 -381 561 -347
rect 729 -381 745 -347
rect 545 -397 745 -381
rect 803 -347 1003 -300
rect 803 -381 819 -347
rect 987 -381 1003 -347
rect 803 -397 1003 -381
<< polycont >>
rect -987 347 -819 381
rect -729 347 -561 381
rect -471 347 -303 381
rect -213 347 -45 381
rect 45 347 213 381
rect 303 347 471 381
rect 561 347 729 381
rect 819 347 987 381
rect -987 -381 -819 -347
rect -729 -381 -561 -347
rect -471 -381 -303 -347
rect -213 -381 -45 -347
rect 45 -381 213 -347
rect 303 -381 471 -347
rect 561 -381 729 -347
rect 819 -381 987 -347
<< locali >>
rect -1183 485 -1087 519
rect 1087 485 1183 519
rect -1183 423 -1149 485
rect 1149 423 1183 485
rect -1003 347 -987 381
rect -819 347 -803 381
rect -745 347 -729 381
rect -561 347 -545 381
rect -487 347 -471 381
rect -303 347 -287 381
rect -229 347 -213 381
rect -45 347 -29 381
rect 29 347 45 381
rect 213 347 229 381
rect 287 347 303 381
rect 471 347 487 381
rect 545 347 561 381
rect 729 347 745 381
rect 803 347 819 381
rect 987 347 1003 381
rect -1049 288 -1015 304
rect -1049 -304 -1015 -288
rect -791 288 -757 304
rect -791 -304 -757 -288
rect -533 288 -499 304
rect -533 -304 -499 -288
rect -275 288 -241 304
rect -275 -304 -241 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 241 288 275 304
rect 241 -304 275 -288
rect 499 288 533 304
rect 499 -304 533 -288
rect 757 288 791 304
rect 757 -304 791 -288
rect 1015 288 1049 304
rect 1015 -304 1049 -288
rect -1003 -381 -987 -347
rect -819 -381 -803 -347
rect -745 -381 -729 -347
rect -561 -381 -545 -347
rect -487 -381 -471 -347
rect -303 -381 -287 -347
rect -229 -381 -213 -347
rect -45 -381 -29 -347
rect 29 -381 45 -347
rect 213 -381 229 -347
rect 287 -381 303 -347
rect 471 -381 487 -347
rect 545 -381 561 -347
rect 729 -381 745 -347
rect 803 -381 819 -347
rect 987 -381 1003 -347
rect 1149 -485 1183 -423
rect -1183 -519 -1087 -485
rect 1087 -519 1183 -485
<< viali >>
rect -987 347 -819 381
rect -729 347 -561 381
rect -471 347 -303 381
rect -213 347 -45 381
rect 45 347 213 381
rect 303 347 471 381
rect 561 347 729 381
rect 819 347 987 381
rect -1183 -423 -1149 0
rect -1049 41 -1015 271
rect -791 -271 -757 -41
rect -533 41 -499 271
rect -275 -271 -241 -41
rect -17 41 17 271
rect 241 -271 275 -41
rect 499 41 533 271
rect 757 -271 791 -41
rect 1015 41 1049 271
rect -987 -381 -819 -347
rect -729 -381 -561 -347
rect -471 -381 -303 -347
rect -213 -381 -45 -347
rect 45 -381 213 -347
rect 303 -381 471 -347
rect 561 -381 729 -347
rect 819 -381 987 -347
rect -1183 -485 -1149 -423
<< metal1 >>
rect -999 381 -807 387
rect -999 347 -987 381
rect -819 347 -807 381
rect -999 341 -807 347
rect -741 381 -549 387
rect -741 347 -729 381
rect -561 347 -549 381
rect -741 341 -549 347
rect -483 381 -291 387
rect -483 347 -471 381
rect -303 347 -291 381
rect -483 341 -291 347
rect -225 381 -33 387
rect -225 347 -213 381
rect -45 347 -33 381
rect -225 341 -33 347
rect 33 381 225 387
rect 33 347 45 381
rect 213 347 225 381
rect 33 341 225 347
rect 291 381 483 387
rect 291 347 303 381
rect 471 347 483 381
rect 291 341 483 347
rect 549 381 741 387
rect 549 347 561 381
rect 729 347 741 381
rect 549 341 741 347
rect 807 381 999 387
rect 807 347 819 381
rect 987 347 999 381
rect 807 341 999 347
rect -1055 271 -1009 283
rect -1055 41 -1049 271
rect -1015 41 -1009 271
rect -1055 29 -1009 41
rect -539 271 -493 283
rect -539 41 -533 271
rect -499 41 -493 271
rect -539 29 -493 41
rect -23 271 23 283
rect -23 41 -17 271
rect 17 41 23 271
rect -23 29 23 41
rect 493 271 539 283
rect 493 41 499 271
rect 533 41 539 271
rect 493 29 539 41
rect 1009 271 1055 283
rect 1009 41 1015 271
rect 1049 41 1055 271
rect 1009 29 1055 41
rect -1189 0 -1143 12
rect -1189 -485 -1183 0
rect -1149 -485 -1143 0
rect -797 -41 -751 -29
rect -797 -271 -791 -41
rect -757 -271 -751 -41
rect -797 -283 -751 -271
rect -281 -41 -235 -29
rect -281 -271 -275 -41
rect -241 -271 -235 -41
rect -281 -283 -235 -271
rect 235 -41 281 -29
rect 235 -271 241 -41
rect 275 -271 281 -41
rect 235 -283 281 -271
rect 751 -41 797 -29
rect 751 -271 757 -41
rect 791 -271 797 -41
rect 751 -283 797 -271
rect -999 -347 -807 -341
rect -999 -381 -987 -347
rect -819 -381 -807 -347
rect -999 -387 -807 -381
rect -741 -347 -549 -341
rect -741 -381 -729 -347
rect -561 -381 -549 -347
rect -741 -387 -549 -381
rect -483 -347 -291 -341
rect -483 -381 -471 -347
rect -303 -381 -291 -347
rect -483 -387 -291 -381
rect -225 -347 -33 -341
rect -225 -381 -213 -347
rect -45 -381 -33 -347
rect -225 -387 -33 -381
rect 33 -347 225 -341
rect 33 -381 45 -347
rect 213 -381 225 -347
rect 33 -387 225 -381
rect 291 -347 483 -341
rect 291 -381 303 -347
rect 471 -381 483 -347
rect 291 -387 483 -381
rect 549 -347 741 -341
rect 549 -381 561 -347
rect 729 -381 741 -347
rect 549 -387 741 -381
rect 807 -347 999 -341
rect 807 -381 819 -347
rect 987 -381 999 -347
rect 807 -387 999 -381
rect -1189 -497 -1143 -485
<< properties >>
string FIXED_BBOX -1166 -502 1166 502
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 3.0 l 1.0 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl +50 viagt 0
<< end >>
