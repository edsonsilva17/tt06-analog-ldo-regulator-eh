magic
tech sky130A
magscale 1 2
timestamp 1713025156
<< metal1 >>
rect 13650 20300 15430 20420
rect 13650 10840 13770 20300
rect 15470 12870 15590 17210
rect 31060 13080 31430 13200
rect 15470 12770 15480 12870
rect 15580 12770 15590 12870
rect 15470 12760 15590 12770
rect 13650 10750 13660 10840
rect 13760 10750 13770 10840
rect 13650 10740 13770 10750
rect 15440 8170 15560 9680
rect 31310 8310 31430 13080
rect 31310 8220 31320 8310
rect 31420 8220 31430 8310
rect 31310 8210 31430 8220
rect 15440 8160 22600 8170
rect 15440 8060 22490 8160
rect 22590 8060 22600 8160
rect 15440 8050 22600 8060
rect 26890 2750 31060 2760
rect 26890 2650 26900 2750
rect 27010 2650 31060 2750
rect 26890 2640 31060 2650
<< via1 >>
rect 15480 12770 15580 12870
rect 13660 10750 13760 10840
rect 31320 8220 31420 8310
rect 22490 8060 22590 8160
rect 26900 2650 27010 2750
<< metal2 >>
rect 15470 12870 15590 12880
rect 15470 12770 15480 12870
rect 15580 12770 15590 12870
rect 13660 10840 13760 10850
rect 13660 10740 13760 10750
rect 15470 7340 15590 12770
rect 31320 8310 31420 8320
rect 31320 8210 31420 8220
rect 22490 8160 22590 8170
rect 22490 8050 22590 8060
rect 15470 7230 15480 7340
rect 15580 7230 15590 7340
rect 15470 7220 15590 7230
rect 26900 2750 27010 2760
rect 26900 2640 27010 2650
<< via2 >>
rect 13660 10750 13760 10840
rect 31320 8220 31420 8310
rect 22490 8060 22590 8160
rect 15480 7230 15580 7340
rect 26900 2650 27010 2750
<< metal3 >>
rect 13650 10840 13770 10845
rect 13650 10750 13660 10840
rect 13760 10750 13770 10840
rect 13650 10745 13770 10750
rect 31310 8310 31430 8315
rect 31310 8220 31320 8310
rect 31420 8220 31430 8310
rect 31310 8215 31430 8220
rect 22480 8160 22600 8165
rect 22480 8060 22490 8160
rect 22590 8060 22600 8160
rect 22480 8055 22600 8060
rect 15470 7340 15590 7345
rect 15470 7230 15480 7340
rect 15580 7230 18180 7340
rect 15470 7220 18180 7230
rect 18060 6950 18180 7220
rect 18060 6850 18070 6950
rect 18170 6850 18180 6950
rect 18060 6840 18180 6850
rect 26890 2750 27020 2755
rect 26890 2650 26900 2750
rect 27010 2650 27020 2750
rect 26890 2645 27020 2650
<< via3 >>
rect 13660 10750 13760 10840
rect 31320 8220 31420 8310
rect 22490 8060 22590 8160
rect 18070 6850 18170 6950
rect 26900 2650 27010 2750
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 1000 500 44152
rect 9800 1000 10100 44152
rect 13648 10840 13768 10852
rect 13648 10750 13660 10840
rect 13760 10750 13768 10840
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 10750
rect 31310 8326 31430 8330
rect 31310 8310 31432 8326
rect 31310 8220 31320 8310
rect 31420 8220 31432 8310
rect 31310 8210 31432 8220
rect 22480 8160 22600 8170
rect 22480 8060 22490 8160
rect 22590 8060 22600 8160
rect 18065 6950 18183 6965
rect 18065 6850 18070 6950
rect 18170 6850 18183 6950
rect 18065 200 18183 6850
rect 18064 0 18184 200
rect 22480 0 22600 8060
rect 26890 2750 27020 2760
rect 26890 2650 26900 2750
rect 27010 2650 27020 2750
rect 26890 2380 27020 2650
rect 26896 0 27016 2380
rect 31312 715 31432 8210
rect 31314 200 31431 715
rect 31312 0 31432 200
use top-1  top-1_0
timestamp 1712983369
transform -1 0 30830 0 -1 29420
box -230 600 15430 26820
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
