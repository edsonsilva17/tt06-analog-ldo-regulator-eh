VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_edsonsilva17_ldo
  CLASS BLOCK ;
  FOREIGN tt_um_edsonsilva17_ldo ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 80.760 81.060 83.540 100.140 ;
      LAYER nwell ;
        RECT 83.820 85.830 86.900 95.400 ;
        RECT 88.940 88.900 101.550 100.150 ;
        RECT 88.940 82.930 108.000 88.900 ;
      LAYER pwell ;
        RECT 88.920 77.060 99.940 82.640 ;
        RECT 82.385 49.815 94.965 52.595 ;
      LAYER nwell ;
        RECT 142.580 46.910 147.450 57.100 ;
        RECT 148.780 54.910 153.650 65.100 ;
      LAYER li1 ;
        RECT 81.000 99.730 83.300 99.900 ;
        RECT 81.000 90.970 81.170 99.730 ;
        RECT 81.900 99.040 82.400 99.210 ;
        RECT 81.670 91.830 81.840 98.870 ;
        RECT 82.460 91.830 82.630 98.870 ;
        RECT 81.900 91.490 82.400 91.660 ;
        RECT 83.130 90.970 83.300 99.730 ;
        RECT 89.330 99.590 101.160 99.760 ;
        RECT 81.000 90.800 83.300 90.970 ;
        RECT 84.210 94.840 86.510 95.010 ;
        RECT 84.210 90.990 84.380 94.840 ;
        RECT 85.110 94.150 85.610 94.320 ;
        RECT 84.880 91.895 85.050 93.935 ;
        RECT 85.670 91.895 85.840 93.935 ;
        RECT 85.110 91.510 85.610 91.680 ;
        RECT 86.340 90.990 86.510 94.840 ;
        RECT 89.330 94.740 89.500 99.590 ;
        RECT 90.230 98.900 91.230 99.070 ;
        RECT 91.520 98.900 92.520 99.070 ;
        RECT 92.810 98.900 93.810 99.070 ;
        RECT 94.100 98.900 95.100 99.070 ;
        RECT 95.390 98.900 96.390 99.070 ;
        RECT 96.680 98.900 97.680 99.070 ;
        RECT 97.970 98.900 98.970 99.070 ;
        RECT 99.260 98.900 100.260 99.070 ;
        RECT 90.000 95.645 90.170 98.685 ;
        RECT 91.290 95.645 91.460 98.685 ;
        RECT 92.580 95.645 92.750 98.685 ;
        RECT 93.870 95.645 94.040 98.685 ;
        RECT 95.160 95.645 95.330 98.685 ;
        RECT 96.450 95.645 96.620 98.685 ;
        RECT 97.740 95.645 97.910 98.685 ;
        RECT 99.030 95.645 99.200 98.685 ;
        RECT 100.320 95.645 100.490 98.685 ;
        RECT 90.230 95.260 91.230 95.430 ;
        RECT 91.520 95.260 92.520 95.430 ;
        RECT 92.810 95.260 93.810 95.430 ;
        RECT 94.100 95.260 95.100 95.430 ;
        RECT 95.390 95.260 96.390 95.430 ;
        RECT 96.680 95.260 97.680 95.430 ;
        RECT 97.970 95.260 98.970 95.430 ;
        RECT 99.260 95.260 100.260 95.430 ;
        RECT 100.990 94.740 101.160 99.590 ;
        RECT 89.330 94.570 101.160 94.740 ;
        RECT 84.210 90.820 86.510 90.990 ;
        RECT 89.330 93.940 101.160 94.110 ;
        RECT 81.000 90.230 83.300 90.400 ;
        RECT 81.000 81.470 81.170 90.230 ;
        RECT 81.900 89.540 82.400 89.710 ;
        RECT 81.670 82.330 81.840 89.370 ;
        RECT 82.460 82.330 82.630 89.370 ;
        RECT 81.900 81.990 82.400 82.160 ;
        RECT 83.130 81.470 83.300 90.230 ;
        RECT 84.210 90.240 86.510 90.410 ;
        RECT 84.210 86.390 84.380 90.240 ;
        RECT 85.110 89.550 85.610 89.720 ;
        RECT 84.880 87.295 85.050 89.335 ;
        RECT 85.670 87.295 85.840 89.335 ;
        RECT 85.110 86.910 85.610 87.080 ;
        RECT 86.340 86.390 86.510 90.240 ;
        RECT 89.330 89.090 89.500 93.940 ;
        RECT 90.230 93.250 91.230 93.420 ;
        RECT 91.520 93.250 92.520 93.420 ;
        RECT 92.810 93.250 93.810 93.420 ;
        RECT 94.100 93.250 95.100 93.420 ;
        RECT 95.390 93.250 96.390 93.420 ;
        RECT 96.680 93.250 97.680 93.420 ;
        RECT 97.970 93.250 98.970 93.420 ;
        RECT 99.260 93.250 100.260 93.420 ;
        RECT 90.000 89.995 90.170 93.035 ;
        RECT 91.290 89.995 91.460 93.035 ;
        RECT 92.580 89.995 92.750 93.035 ;
        RECT 93.870 89.995 94.040 93.035 ;
        RECT 95.160 89.995 95.330 93.035 ;
        RECT 96.450 89.995 96.620 93.035 ;
        RECT 97.740 89.995 97.910 93.035 ;
        RECT 99.030 89.995 99.200 93.035 ;
        RECT 100.320 89.995 100.490 93.035 ;
        RECT 90.230 89.610 91.230 89.780 ;
        RECT 91.520 89.610 92.520 89.780 ;
        RECT 92.810 89.610 93.810 89.780 ;
        RECT 94.100 89.610 95.100 89.780 ;
        RECT 95.390 89.610 96.390 89.780 ;
        RECT 96.680 89.610 97.680 89.780 ;
        RECT 97.970 89.610 98.970 89.780 ;
        RECT 99.260 89.610 100.260 89.780 ;
        RECT 100.990 89.090 101.160 93.940 ;
        RECT 89.330 88.920 101.160 89.090 ;
        RECT 84.210 86.220 86.510 86.390 ;
        RECT 89.330 88.340 107.610 88.510 ;
        RECT 89.330 83.490 89.500 88.340 ;
        RECT 90.230 87.650 91.230 87.820 ;
        RECT 91.520 87.650 92.520 87.820 ;
        RECT 92.810 87.650 93.810 87.820 ;
        RECT 94.100 87.650 95.100 87.820 ;
        RECT 95.390 87.650 96.390 87.820 ;
        RECT 96.680 87.650 97.680 87.820 ;
        RECT 97.970 87.650 98.970 87.820 ;
        RECT 99.260 87.650 100.260 87.820 ;
        RECT 100.550 87.650 101.550 87.820 ;
        RECT 101.840 87.650 102.840 87.820 ;
        RECT 103.130 87.650 104.130 87.820 ;
        RECT 104.420 87.650 105.420 87.820 ;
        RECT 105.710 87.650 106.710 87.820 ;
        RECT 90.000 84.395 90.170 87.435 ;
        RECT 91.290 84.395 91.460 87.435 ;
        RECT 92.580 84.395 92.750 87.435 ;
        RECT 93.870 84.395 94.040 87.435 ;
        RECT 95.160 84.395 95.330 87.435 ;
        RECT 96.450 84.395 96.620 87.435 ;
        RECT 97.740 84.395 97.910 87.435 ;
        RECT 99.030 84.395 99.200 87.435 ;
        RECT 100.320 84.395 100.490 87.435 ;
        RECT 101.610 84.395 101.780 87.435 ;
        RECT 102.900 84.395 103.070 87.435 ;
        RECT 104.190 84.395 104.360 87.435 ;
        RECT 105.480 84.395 105.650 87.435 ;
        RECT 106.770 84.395 106.940 87.435 ;
        RECT 90.230 84.010 91.230 84.180 ;
        RECT 91.520 84.010 92.520 84.180 ;
        RECT 92.810 84.010 93.810 84.180 ;
        RECT 94.100 84.010 95.100 84.180 ;
        RECT 95.390 84.010 96.390 84.180 ;
        RECT 96.680 84.010 97.680 84.180 ;
        RECT 97.970 84.010 98.970 84.180 ;
        RECT 99.260 84.010 100.260 84.180 ;
        RECT 100.550 84.010 101.550 84.180 ;
        RECT 101.840 84.010 102.840 84.180 ;
        RECT 103.130 84.010 104.130 84.180 ;
        RECT 104.420 84.010 105.420 84.180 ;
        RECT 105.710 84.010 106.710 84.180 ;
        RECT 107.440 83.490 107.610 88.340 ;
        RECT 89.330 83.320 107.610 83.490 ;
        RECT 81.000 81.300 83.300 81.470 ;
        RECT 89.160 82.230 99.700 82.400 ;
        RECT 89.160 77.470 89.330 82.230 ;
        RECT 90.060 81.540 91.060 81.710 ;
        RECT 91.350 81.540 92.350 81.710 ;
        RECT 92.640 81.540 93.640 81.710 ;
        RECT 93.930 81.540 94.930 81.710 ;
        RECT 95.220 81.540 96.220 81.710 ;
        RECT 96.510 81.540 97.510 81.710 ;
        RECT 97.800 81.540 98.800 81.710 ;
        RECT 89.830 78.330 90.000 81.370 ;
        RECT 91.120 78.330 91.290 81.370 ;
        RECT 92.410 78.330 92.580 81.370 ;
        RECT 93.700 78.330 93.870 81.370 ;
        RECT 94.990 78.330 95.160 81.370 ;
        RECT 96.280 78.330 96.450 81.370 ;
        RECT 97.570 78.330 97.740 81.370 ;
        RECT 98.860 78.330 99.030 81.370 ;
        RECT 90.060 77.990 91.060 78.160 ;
        RECT 91.350 77.990 92.350 78.160 ;
        RECT 92.640 77.990 93.640 78.160 ;
        RECT 93.930 77.990 94.930 78.160 ;
        RECT 95.220 77.990 96.220 78.160 ;
        RECT 96.510 77.990 97.510 78.160 ;
        RECT 97.800 77.990 98.800 78.160 ;
        RECT 99.530 77.470 99.700 82.230 ;
        RECT 89.160 77.300 99.700 77.470 ;
        RECT 148.960 64.750 153.470 64.920 ;
        RECT 142.760 56.750 147.270 56.920 ;
        RECT 82.625 52.185 94.725 52.355 ;
        RECT 82.625 50.225 82.795 52.185 ;
        RECT 83.655 51.515 93.695 51.685 ;
        RECT 83.315 50.955 83.485 51.455 ;
        RECT 93.865 50.955 94.035 51.455 ;
        RECT 83.655 50.725 93.695 50.895 ;
        RECT 94.555 50.225 94.725 52.185 ;
        RECT 82.625 50.055 94.725 50.225 ;
        RECT 142.760 47.260 142.930 56.750 ;
        RECT 143.560 56.240 143.910 56.410 ;
        RECT 144.200 56.240 144.550 56.410 ;
        RECT 144.840 56.240 145.190 56.410 ;
        RECT 145.480 56.240 145.830 56.410 ;
        RECT 146.120 56.240 146.470 56.410 ;
        RECT 143.330 47.985 143.500 56.025 ;
        RECT 143.970 47.985 144.140 56.025 ;
        RECT 144.610 47.985 144.780 56.025 ;
        RECT 145.250 47.985 145.420 56.025 ;
        RECT 145.890 47.985 146.060 56.025 ;
        RECT 146.530 47.985 146.700 56.025 ;
        RECT 143.560 47.600 143.910 47.770 ;
        RECT 144.200 47.600 144.550 47.770 ;
        RECT 144.840 47.600 145.190 47.770 ;
        RECT 145.480 47.600 145.830 47.770 ;
        RECT 146.120 47.600 146.470 47.770 ;
        RECT 147.100 47.260 147.270 56.750 ;
        RECT 148.960 55.260 149.130 64.750 ;
        RECT 149.760 64.240 150.110 64.410 ;
        RECT 150.400 64.240 150.750 64.410 ;
        RECT 151.040 64.240 151.390 64.410 ;
        RECT 151.680 64.240 152.030 64.410 ;
        RECT 152.320 64.240 152.670 64.410 ;
        RECT 149.530 55.985 149.700 64.025 ;
        RECT 150.170 55.985 150.340 64.025 ;
        RECT 150.810 55.985 150.980 64.025 ;
        RECT 151.450 55.985 151.620 64.025 ;
        RECT 152.090 55.985 152.260 64.025 ;
        RECT 152.730 55.985 152.900 64.025 ;
        RECT 149.760 55.600 150.110 55.770 ;
        RECT 150.400 55.600 150.750 55.770 ;
        RECT 151.040 55.600 151.390 55.770 ;
        RECT 151.680 55.600 152.030 55.770 ;
        RECT 152.320 55.600 152.670 55.770 ;
        RECT 153.300 55.260 153.470 64.750 ;
        RECT 148.960 55.090 153.470 55.260 ;
        RECT 142.760 47.090 147.270 47.260 ;
      LAYER mcon ;
        RECT 81.980 99.040 82.320 99.210 ;
        RECT 81.670 91.995 81.840 94.060 ;
        RECT 82.460 91.995 82.630 94.060 ;
        RECT 81.980 91.490 82.320 91.660 ;
        RECT 85.190 94.150 85.530 94.320 ;
        RECT 84.880 91.975 85.050 93.855 ;
        RECT 85.670 91.975 85.840 93.855 ;
        RECT 90.310 98.900 91.150 99.070 ;
        RECT 91.600 98.900 92.440 99.070 ;
        RECT 92.890 98.900 93.730 99.070 ;
        RECT 94.180 98.900 95.020 99.070 ;
        RECT 95.470 98.900 96.310 99.070 ;
        RECT 96.760 98.900 97.600 99.070 ;
        RECT 98.050 98.900 98.890 99.070 ;
        RECT 99.340 98.900 100.180 99.070 ;
        RECT 90.000 95.810 90.170 96.960 ;
        RECT 91.290 97.370 91.460 98.520 ;
        RECT 92.580 95.810 92.750 96.960 ;
        RECT 93.870 97.370 94.040 98.520 ;
        RECT 95.160 95.810 95.330 96.960 ;
        RECT 96.450 97.370 96.620 98.520 ;
        RECT 97.740 95.810 97.910 96.960 ;
        RECT 99.030 97.370 99.200 98.520 ;
        RECT 100.320 95.810 100.490 96.960 ;
        RECT 90.310 95.260 91.150 95.430 ;
        RECT 91.600 95.260 92.440 95.430 ;
        RECT 92.890 95.260 93.730 95.430 ;
        RECT 94.180 95.260 95.020 95.430 ;
        RECT 95.470 95.260 96.310 95.430 ;
        RECT 96.760 95.260 97.600 95.430 ;
        RECT 98.050 95.260 98.890 95.430 ;
        RECT 99.340 95.260 100.180 95.430 ;
        RECT 86.340 92.625 86.510 93.205 ;
        RECT 85.190 91.510 85.530 91.680 ;
        RECT 81.000 87.600 81.170 90.230 ;
        RECT 81.980 89.540 82.320 89.710 ;
        RECT 81.670 87.140 81.840 89.205 ;
        RECT 82.460 87.140 82.630 89.205 ;
        RECT 81.980 81.990 82.320 82.160 ;
        RECT 85.190 89.550 85.530 89.720 ;
        RECT 84.880 87.375 85.050 89.255 ;
        RECT 85.670 87.375 85.840 89.255 ;
        RECT 90.310 93.250 91.150 93.420 ;
        RECT 91.600 93.250 92.440 93.420 ;
        RECT 92.890 93.250 93.730 93.420 ;
        RECT 94.180 93.250 95.020 93.420 ;
        RECT 95.470 93.250 96.310 93.420 ;
        RECT 96.760 93.250 97.600 93.420 ;
        RECT 98.050 93.250 98.890 93.420 ;
        RECT 99.340 93.250 100.180 93.420 ;
        RECT 90.000 90.160 90.170 91.310 ;
        RECT 91.290 91.720 91.460 92.870 ;
        RECT 92.580 90.160 92.750 91.310 ;
        RECT 93.870 91.720 94.040 92.870 ;
        RECT 95.160 90.160 95.330 91.310 ;
        RECT 96.450 91.720 96.620 92.870 ;
        RECT 97.740 90.160 97.910 91.310 ;
        RECT 99.030 91.720 99.200 92.870 ;
        RECT 100.320 90.160 100.490 91.310 ;
        RECT 100.990 91.515 101.160 93.940 ;
        RECT 90.310 89.610 91.150 89.780 ;
        RECT 91.600 89.610 92.440 89.780 ;
        RECT 92.890 89.610 93.730 89.780 ;
        RECT 94.180 89.610 95.020 89.780 ;
        RECT 95.470 89.610 96.310 89.780 ;
        RECT 96.760 89.610 97.600 89.780 ;
        RECT 98.050 89.610 98.890 89.780 ;
        RECT 99.340 89.610 100.180 89.780 ;
        RECT 86.340 88.025 86.510 88.605 ;
        RECT 85.190 86.910 85.530 87.080 ;
        RECT 90.310 87.650 91.150 87.820 ;
        RECT 91.600 87.650 92.440 87.820 ;
        RECT 92.890 87.650 93.730 87.820 ;
        RECT 94.180 87.650 95.020 87.820 ;
        RECT 95.470 87.650 96.310 87.820 ;
        RECT 96.760 87.650 97.600 87.820 ;
        RECT 98.050 87.650 98.890 87.820 ;
        RECT 99.340 87.650 100.180 87.820 ;
        RECT 100.630 87.650 101.470 87.820 ;
        RECT 101.920 87.650 102.760 87.820 ;
        RECT 103.210 87.650 104.050 87.820 ;
        RECT 104.500 87.650 105.340 87.820 ;
        RECT 105.790 87.650 106.630 87.820 ;
        RECT 90.000 86.120 90.170 87.270 ;
        RECT 91.290 84.560 91.460 85.710 ;
        RECT 92.580 86.120 92.750 87.270 ;
        RECT 93.870 84.560 94.040 85.710 ;
        RECT 95.160 86.120 95.330 87.270 ;
        RECT 96.450 84.560 96.620 85.710 ;
        RECT 97.740 86.120 97.910 87.270 ;
        RECT 99.030 84.560 99.200 85.710 ;
        RECT 100.320 86.120 100.490 87.270 ;
        RECT 101.610 84.560 101.780 85.710 ;
        RECT 102.900 86.120 103.070 87.270 ;
        RECT 104.190 84.560 104.360 85.710 ;
        RECT 105.480 86.120 105.650 87.270 ;
        RECT 106.770 84.560 106.940 85.710 ;
        RECT 107.440 85.915 107.610 88.340 ;
        RECT 90.310 84.010 91.150 84.180 ;
        RECT 91.600 84.010 92.440 84.180 ;
        RECT 92.890 84.010 93.730 84.180 ;
        RECT 94.180 84.010 95.020 84.180 ;
        RECT 95.470 84.010 96.310 84.180 ;
        RECT 96.760 84.010 97.600 84.180 ;
        RECT 98.050 84.010 98.890 84.180 ;
        RECT 99.340 84.010 100.180 84.180 ;
        RECT 100.630 84.010 101.470 84.180 ;
        RECT 101.920 84.010 102.760 84.180 ;
        RECT 103.210 84.010 104.050 84.180 ;
        RECT 104.500 84.010 105.340 84.180 ;
        RECT 105.790 84.010 106.630 84.180 ;
        RECT 90.140 81.540 90.980 81.710 ;
        RECT 91.430 81.540 92.270 81.710 ;
        RECT 92.720 81.540 93.560 81.710 ;
        RECT 94.010 81.540 94.850 81.710 ;
        RECT 95.300 81.540 96.140 81.710 ;
        RECT 96.590 81.540 97.430 81.710 ;
        RECT 97.880 81.540 98.720 81.710 ;
        RECT 89.830 80.055 90.000 81.205 ;
        RECT 91.120 78.495 91.290 79.645 ;
        RECT 92.410 80.055 92.580 81.205 ;
        RECT 93.700 78.495 93.870 79.645 ;
        RECT 94.990 80.055 95.160 81.205 ;
        RECT 96.280 78.495 96.450 79.645 ;
        RECT 97.570 80.055 97.740 81.205 ;
        RECT 98.860 78.495 99.030 79.645 ;
        RECT 99.530 79.850 99.700 82.230 ;
        RECT 90.140 77.990 90.980 78.160 ;
        RECT 91.430 77.990 92.270 78.160 ;
        RECT 92.720 77.990 93.560 78.160 ;
        RECT 94.010 77.990 94.850 78.160 ;
        RECT 95.300 77.990 96.140 78.160 ;
        RECT 96.590 77.990 97.430 78.160 ;
        RECT 97.880 77.990 98.720 78.160 ;
        RECT 87.795 52.185 89.555 52.355 ;
        RECT 91.555 51.515 93.530 51.685 ;
        RECT 83.315 51.035 83.485 51.375 ;
        RECT 93.865 51.035 94.035 51.375 ;
        RECT 83.820 50.725 85.795 50.895 ;
        RECT 143.640 56.240 143.830 56.410 ;
        RECT 144.280 56.240 144.470 56.410 ;
        RECT 144.920 56.240 145.110 56.410 ;
        RECT 145.560 56.240 145.750 56.410 ;
        RECT 146.200 56.240 146.390 56.410 ;
        RECT 143.330 52.710 143.500 55.860 ;
        RECT 143.970 48.150 144.140 51.300 ;
        RECT 144.610 52.710 144.780 55.860 ;
        RECT 145.250 48.150 145.420 51.300 ;
        RECT 145.890 52.710 146.060 55.860 ;
        RECT 146.530 48.150 146.700 51.300 ;
        RECT 143.640 47.600 143.830 47.770 ;
        RECT 144.280 47.600 144.470 47.770 ;
        RECT 144.920 47.600 145.110 47.770 ;
        RECT 145.560 47.600 145.750 47.770 ;
        RECT 146.200 47.600 146.390 47.770 ;
        RECT 149.840 64.240 150.030 64.410 ;
        RECT 150.480 64.240 150.670 64.410 ;
        RECT 151.120 64.240 151.310 64.410 ;
        RECT 151.760 64.240 151.950 64.410 ;
        RECT 152.400 64.240 152.590 64.410 ;
        RECT 149.530 60.710 149.700 63.860 ;
        RECT 150.170 56.150 150.340 59.300 ;
        RECT 150.810 60.710 150.980 63.860 ;
        RECT 151.450 56.150 151.620 59.300 ;
        RECT 152.090 60.710 152.260 63.860 ;
        RECT 152.730 56.150 152.900 59.300 ;
        RECT 149.840 55.600 150.030 55.770 ;
        RECT 150.480 55.600 150.670 55.770 ;
        RECT 151.120 55.600 151.310 55.770 ;
        RECT 151.760 55.600 151.950 55.770 ;
        RECT 152.400 55.600 152.590 55.770 ;
        RECT 150.175 55.090 152.255 55.260 ;
        RECT 143.975 47.090 146.055 47.260 ;
      LAYER met1 ;
        RECT 76.400 102.200 77.400 102.300 ;
        RECT 76.400 102.100 108.400 102.200 ;
        RECT 68.250 101.500 108.400 102.100 ;
        RECT 68.250 53.700 68.850 101.500 ;
        RECT 76.400 101.400 108.400 101.500 ;
        RECT 76.400 101.300 77.400 101.400 ;
        RECT 107.600 100.650 108.400 101.400 ;
        RECT 107.500 99.650 108.500 100.650 ;
        RECT 81.920 99.010 82.380 99.240 ;
        RECT 90.200 98.750 102.450 99.200 ;
        RECT 91.260 98.300 91.490 98.580 ;
        RECT 93.840 98.300 94.070 98.580 ;
        RECT 96.420 98.300 96.650 98.580 ;
        RECT 99.000 98.300 99.230 98.580 ;
        RECT 102.000 98.300 102.450 98.750 ;
        RECT 107.600 98.400 108.400 99.650 ;
        RECT 107.500 98.300 108.500 98.400 ;
        RECT 91.250 97.550 108.500 98.300 ;
        RECT 91.260 97.310 91.490 97.550 ;
        RECT 93.840 97.310 94.070 97.550 ;
        RECT 96.420 97.310 96.650 97.550 ;
        RECT 99.000 97.310 99.230 97.550 ;
        RECT 107.500 97.400 108.500 97.550 ;
        RECT 89.970 96.750 90.200 97.020 ;
        RECT 92.550 96.750 92.780 97.020 ;
        RECT 95.130 96.750 95.360 97.020 ;
        RECT 97.710 96.750 97.940 97.020 ;
        RECT 100.290 96.750 100.520 97.020 ;
        RECT 100.960 96.750 101.190 97.225 ;
        RECT 79.800 95.900 80.800 96.150 ;
        RECT 89.970 96.000 108.400 96.750 ;
        RECT 79.800 95.400 85.600 95.900 ;
        RECT 89.970 95.750 90.200 96.000 ;
        RECT 92.550 95.750 92.780 96.000 ;
        RECT 95.130 95.750 95.360 96.000 ;
        RECT 97.710 95.750 97.940 96.000 ;
        RECT 100.290 95.750 100.520 96.000 ;
        RECT 79.800 95.150 80.800 95.400 ;
        RECT 79.900 94.400 80.700 95.150 ;
        RECT 80.970 93.300 81.200 93.660 ;
        RECT 81.640 93.300 81.870 94.120 ;
        RECT 79.900 92.550 81.870 93.300 ;
        RECT 79.900 91.100 80.700 92.550 ;
        RECT 77.550 91.000 78.550 91.100 ;
        RECT 79.800 91.000 80.800 91.100 ;
        RECT 77.550 90.200 80.800 91.000 ;
        RECT 80.970 90.910 81.200 92.550 ;
        RECT 81.640 91.935 81.870 92.550 ;
        RECT 82.430 93.300 82.660 94.120 ;
        RECT 85.100 94.100 85.600 95.400 ;
        RECT 90.250 95.230 91.210 95.460 ;
        RECT 91.540 95.230 92.500 95.460 ;
        RECT 92.830 95.230 93.790 95.460 ;
        RECT 94.120 95.230 95.080 95.460 ;
        RECT 95.410 95.230 96.370 95.460 ;
        RECT 96.700 95.230 97.660 95.460 ;
        RECT 97.990 95.230 98.950 95.460 ;
        RECT 99.280 95.230 100.240 95.460 ;
        RECT 100.960 94.680 101.190 96.000 ;
        RECT 84.850 93.300 85.080 93.915 ;
        RECT 82.430 92.550 85.080 93.300 ;
        RECT 82.430 91.935 82.660 92.550 ;
        RECT 81.900 90.750 82.400 91.700 ;
        RECT 83.400 90.750 83.900 92.550 ;
        RECT 84.850 91.915 85.080 92.550 ;
        RECT 85.640 93.300 85.870 93.915 ;
        RECT 85.640 92.550 87.750 93.300 ;
        RECT 90.250 93.220 91.210 93.450 ;
        RECT 91.540 93.220 92.500 93.450 ;
        RECT 92.830 93.220 93.790 93.450 ;
        RECT 94.120 93.220 95.080 93.450 ;
        RECT 95.410 93.220 96.370 93.450 ;
        RECT 96.700 93.220 97.660 93.450 ;
        RECT 97.990 93.220 98.950 93.450 ;
        RECT 99.280 93.220 100.240 93.450 ;
        RECT 85.640 91.915 85.870 92.550 ;
        RECT 85.130 91.480 85.590 91.710 ;
        RECT 81.900 90.450 83.900 90.750 ;
        RECT 86.600 91.100 87.750 92.550 ;
        RECT 91.260 92.650 91.490 92.930 ;
        RECT 93.840 92.650 94.070 92.930 ;
        RECT 96.420 92.650 96.650 92.930 ;
        RECT 99.000 92.650 99.230 92.930 ;
        RECT 100.960 92.650 101.190 94.000 ;
        RECT 107.600 92.750 108.400 96.000 ;
        RECT 107.500 92.650 108.500 92.750 ;
        RECT 91.260 91.900 108.500 92.650 ;
        RECT 91.260 91.660 91.490 91.900 ;
        RECT 93.840 91.660 94.070 91.900 ;
        RECT 96.420 91.660 96.650 91.900 ;
        RECT 99.000 91.660 99.230 91.900 ;
        RECT 100.960 91.455 101.190 91.900 ;
        RECT 107.500 91.750 108.500 91.900 ;
        RECT 89.970 91.100 90.200 91.370 ;
        RECT 92.550 91.100 92.780 91.370 ;
        RECT 95.130 91.100 95.360 91.370 ;
        RECT 97.710 91.100 97.940 91.370 ;
        RECT 100.290 91.100 100.520 91.370 ;
        RECT 77.550 90.100 78.550 90.200 ;
        RECT 78.750 87.950 79.550 90.200 ;
        RECT 79.800 90.100 80.800 90.200 ;
        RECT 79.900 88.700 80.700 90.100 ;
        RECT 80.970 88.700 81.200 90.290 ;
        RECT 81.900 89.500 82.400 90.450 ;
        RECT 86.600 90.350 100.520 91.100 ;
        RECT 85.130 89.520 85.590 89.750 ;
        RECT 81.640 88.700 81.870 89.265 ;
        RECT 79.900 87.950 81.870 88.700 ;
        RECT 80.970 87.540 81.200 87.950 ;
        RECT 81.640 87.080 81.870 87.950 ;
        RECT 82.430 88.700 82.660 89.265 ;
        RECT 84.850 88.700 85.080 89.315 ;
        RECT 82.430 87.950 85.080 88.700 ;
        RECT 82.430 87.080 82.660 87.950 ;
        RECT 84.850 87.315 85.080 87.950 ;
        RECT 85.640 88.700 85.870 89.315 ;
        RECT 86.600 88.700 87.750 90.350 ;
        RECT 89.970 90.100 90.200 90.350 ;
        RECT 92.550 90.100 92.780 90.350 ;
        RECT 95.130 90.100 95.360 90.350 ;
        RECT 97.710 90.100 97.940 90.350 ;
        RECT 100.290 90.100 100.520 90.350 ;
        RECT 90.200 89.450 102.450 89.900 ;
        RECT 85.640 87.950 87.750 88.700 ;
        RECT 102.000 88.000 102.450 89.450 ;
        RECT 107.600 88.400 108.400 91.750 ;
        RECT 85.640 87.315 85.870 87.950 ;
        RECT 90.200 87.550 106.700 88.000 ;
        RECT 85.130 87.100 85.590 87.110 ;
        RECT 89.970 87.100 90.200 87.330 ;
        RECT 92.550 87.100 92.780 87.330 ;
        RECT 95.130 87.100 95.360 87.330 ;
        RECT 97.710 87.100 97.940 87.330 ;
        RECT 100.290 87.100 100.520 87.330 ;
        RECT 102.870 87.100 103.100 87.330 ;
        RECT 105.450 87.100 105.680 87.330 ;
        RECT 107.410 87.100 108.400 88.400 ;
        RECT 76.400 85.950 78.550 86.050 ;
        RECT 79.800 85.950 80.800 86.050 ;
        RECT 76.400 85.800 80.800 85.950 ;
        RECT 85.100 85.800 85.600 87.100 ;
        RECT 89.950 86.350 108.400 87.100 ;
        RECT 89.970 86.060 90.200 86.350 ;
        RECT 92.550 86.060 92.780 86.350 ;
        RECT 95.130 86.060 95.360 86.350 ;
        RECT 97.710 86.060 97.940 86.350 ;
        RECT 100.290 86.060 100.520 86.350 ;
        RECT 102.870 86.060 103.100 86.350 ;
        RECT 105.450 86.060 105.680 86.350 ;
        RECT 107.410 85.855 107.640 86.350 ;
        RECT 76.400 85.300 85.600 85.800 ;
        RECT 91.260 85.500 91.490 85.770 ;
        RECT 93.840 85.500 94.070 85.770 ;
        RECT 96.420 85.500 96.650 85.770 ;
        RECT 99.000 85.500 99.230 85.770 ;
        RECT 101.580 85.500 101.810 85.770 ;
        RECT 104.160 85.500 104.390 85.770 ;
        RECT 106.740 85.500 106.970 85.770 ;
        RECT 76.400 85.150 80.800 85.300 ;
        RECT 76.400 85.050 78.550 85.150 ;
        RECT 79.800 85.050 80.800 85.150 ;
        RECT 76.600 63.800 77.200 85.050 ;
        RECT 91.250 84.750 108.400 85.500 ;
        RECT 91.260 84.500 91.490 84.750 ;
        RECT 93.840 84.500 94.070 84.750 ;
        RECT 96.420 84.500 96.650 84.750 ;
        RECT 99.000 84.500 99.230 84.750 ;
        RECT 101.580 84.500 101.810 84.750 ;
        RECT 104.160 84.500 104.390 84.750 ;
        RECT 106.740 84.500 106.970 84.750 ;
        RECT 90.250 83.980 91.210 84.210 ;
        RECT 91.540 83.980 92.500 84.210 ;
        RECT 92.830 83.980 93.790 84.210 ;
        RECT 94.120 83.980 95.080 84.210 ;
        RECT 95.410 83.980 96.370 84.210 ;
        RECT 96.700 83.980 97.660 84.210 ;
        RECT 97.990 83.980 98.950 84.210 ;
        RECT 99.280 83.980 100.240 84.210 ;
        RECT 100.570 83.980 101.530 84.210 ;
        RECT 101.860 83.980 102.820 84.210 ;
        RECT 103.150 83.980 104.110 84.210 ;
        RECT 104.440 83.980 105.400 84.210 ;
        RECT 105.730 83.980 106.690 84.210 ;
        RECT 81.920 81.960 82.380 82.190 ;
        RECT 85.550 81.850 86.100 81.900 ;
        RECT 85.550 81.500 98.800 81.850 ;
        RECT 85.550 81.450 86.100 81.500 ;
        RECT 89.800 81.000 90.030 81.265 ;
        RECT 92.380 81.000 92.610 81.265 ;
        RECT 94.960 81.000 95.190 81.265 ;
        RECT 97.540 81.000 97.770 81.265 ;
        RECT 99.500 81.000 99.730 82.290 ;
        RECT 79.900 80.250 99.750 81.000 ;
        RECT 89.800 79.995 90.030 80.250 ;
        RECT 92.380 79.995 92.610 80.250 ;
        RECT 94.960 79.995 95.190 80.250 ;
        RECT 97.540 79.995 97.770 80.250 ;
        RECT 99.500 79.790 99.730 80.250 ;
        RECT 79.800 79.450 80.800 79.550 ;
        RECT 91.090 79.450 91.320 79.705 ;
        RECT 93.670 79.450 93.900 79.705 ;
        RECT 96.250 79.450 96.480 79.705 ;
        RECT 98.830 79.450 99.060 79.705 ;
        RECT 107.600 79.450 108.400 84.750 ;
        RECT 79.800 78.700 108.400 79.450 ;
        RECT 79.800 78.550 80.800 78.700 ;
        RECT 79.900 51.450 80.700 78.550 ;
        RECT 91.090 78.435 91.320 78.700 ;
        RECT 93.670 78.435 93.900 78.700 ;
        RECT 96.250 78.435 96.480 78.700 ;
        RECT 98.830 78.435 99.060 78.700 ;
        RECT 90.080 77.960 91.040 78.190 ;
        RECT 91.370 77.960 92.330 78.190 ;
        RECT 92.660 77.960 93.620 78.190 ;
        RECT 93.950 77.960 94.910 78.190 ;
        RECT 95.240 77.960 96.200 78.190 ;
        RECT 96.530 77.960 97.490 78.190 ;
        RECT 97.820 77.960 98.780 78.190 ;
        RECT 106.400 66.000 155.300 66.200 ;
        RECT 106.400 65.400 157.150 66.000 ;
        RECT 106.400 65.200 155.300 65.400 ;
        RECT 88.350 52.385 89.000 53.100 ;
        RECT 87.735 52.155 89.615 52.385 ;
        RECT 88.350 52.150 89.000 52.155 ;
        RECT 91.495 51.485 93.590 51.715 ;
        RECT 79.900 51.435 83.500 51.450 ;
        RECT 79.900 50.975 83.515 51.435 ;
        RECT 79.900 50.950 83.500 50.975 ;
        RECT 84.450 50.925 85.200 50.950 ;
        RECT 83.760 50.695 85.855 50.925 ;
        RECT 76.250 49.300 78.400 49.400 ;
        RECT 84.450 49.300 85.200 50.695 ;
        RECT 76.250 48.500 85.200 49.300 ;
        RECT 92.300 49.300 93.050 51.485 ;
        RECT 93.835 50.975 94.065 51.435 ;
        RECT 107.600 49.400 108.400 64.550 ;
        RECT 148.250 63.400 149.250 65.200 ;
        RECT 149.750 64.200 152.750 64.500 ;
        RECT 149.500 63.400 149.730 63.920 ;
        RECT 150.780 63.400 151.010 63.920 ;
        RECT 152.060 63.400 152.290 63.920 ;
        RECT 148.250 62.400 152.350 63.400 ;
        RECT 149.500 60.650 149.730 62.400 ;
        RECT 150.780 60.650 151.010 62.400 ;
        RECT 152.060 60.650 152.290 62.400 ;
        RECT 150.140 59.300 150.370 59.360 ;
        RECT 151.420 59.300 151.650 59.360 ;
        RECT 152.700 59.300 152.930 59.360 ;
        RECT 143.550 56.200 146.450 56.500 ;
        RECT 143.300 54.900 143.530 55.920 ;
        RECT 144.580 54.900 144.810 55.920 ;
        RECT 145.860 54.900 146.090 55.920 ;
        RECT 149.450 55.500 152.950 59.300 ;
        RECT 150.050 54.900 152.350 55.500 ;
        RECT 143.250 53.900 151.650 54.900 ;
        RECT 143.300 52.650 143.530 53.900 ;
        RECT 144.580 52.650 144.810 53.900 ;
        RECT 145.860 52.650 146.090 53.900 ;
        RECT 143.250 49.400 146.750 51.400 ;
        RECT 107.500 49.300 109.650 49.400 ;
        RECT 92.300 48.600 110.950 49.300 ;
        RECT 92.300 48.500 109.650 48.600 ;
        RECT 76.250 48.400 78.400 48.500 ;
        RECT 107.500 48.400 109.650 48.500 ;
        RECT 137.650 48.400 146.750 49.400 ;
        RECT 150.450 49.200 151.250 53.900 ;
        RECT 76.450 40.850 77.050 48.400 ;
        RECT 143.250 47.500 146.750 48.400 ;
        RECT 143.850 46.900 146.150 47.500 ;
        RECT 156.550 41.050 157.150 65.400 ;
        RECT 76.450 40.250 113.000 40.850 ;
        RECT 153.150 14.000 154.150 14.900 ;
        RECT 153.150 13.800 155.300 14.000 ;
        RECT 134.450 13.200 155.300 13.800 ;
        RECT 153.150 13.000 155.300 13.200 ;
      LAYER via ;
        RECT 102.000 97.700 102.450 98.150 ;
        RECT 80.000 94.500 80.600 95.050 ;
        RECT 78.850 88.050 79.450 88.600 ;
        RECT 80.000 88.050 80.600 88.600 ;
        RECT 83.350 88.050 83.900 88.600 ;
        RECT 102.050 89.500 102.400 89.850 ;
        RECT 107.700 89.650 108.300 90.250 ;
        RECT 85.600 81.450 86.050 81.900 ;
        RECT 80.000 80.350 80.600 80.900 ;
        RECT 81.900 78.750 82.300 79.400 ;
        RECT 76.650 63.850 77.150 64.350 ;
        RECT 68.300 53.750 68.800 54.200 ;
        RECT 106.500 65.300 107.300 66.100 ;
        RECT 143.150 65.250 144.050 66.150 ;
        RECT 107.700 63.850 108.300 64.450 ;
        RECT 88.450 52.550 88.900 53.000 ;
        RECT 80.000 48.600 80.600 49.200 ;
        RECT 110.250 48.700 110.850 49.200 ;
        RECT 137.750 48.500 138.550 49.300 ;
        RECT 150.550 49.300 151.150 49.900 ;
        RECT 156.600 41.100 157.100 41.550 ;
        RECT 112.450 40.300 112.950 40.800 ;
        RECT 153.350 14.100 153.950 14.700 ;
        RECT 134.500 13.250 135.050 13.750 ;
      LAYER met2 ;
        RECT 80.000 94.450 80.600 95.100 ;
        RECT 102.000 89.450 102.450 98.200 ;
        RECT 78.750 66.200 79.550 88.700 ;
        RECT 79.900 80.250 80.700 88.700 ;
        RECT 83.350 85.050 83.900 88.650 ;
        RECT 83.350 84.500 86.100 85.050 ;
        RECT 85.550 81.400 86.100 84.500 ;
        RECT 81.900 78.700 82.300 79.450 ;
        RECT 78.750 65.200 107.400 66.200 ;
        RECT 68.300 53.700 68.800 54.250 ;
        RECT 76.600 36.100 77.200 64.400 ;
        RECT 78.750 53.100 79.550 65.200 ;
        RECT 107.600 63.750 108.400 90.300 ;
        RECT 143.150 65.200 144.050 66.200 ;
        RECT 78.750 52.500 89.000 53.100 ;
        RECT 78.750 52.450 88.350 52.500 ;
        RECT 80.000 48.550 80.600 49.250 ;
        RECT 110.250 48.650 110.850 49.250 ;
        RECT 137.750 48.450 138.550 49.350 ;
        RECT 150.550 49.250 151.150 49.950 ;
        RECT 156.600 41.050 157.100 41.600 ;
        RECT 112.450 40.250 112.950 40.850 ;
        RECT 153.350 14.050 153.950 14.750 ;
        RECT 134.500 13.200 135.050 13.800 ;
      LAYER via2 ;
        RECT 80.000 94.500 80.600 95.050 ;
        RECT 85.600 81.450 86.050 81.900 ;
        RECT 81.900 78.750 82.300 79.400 ;
        RECT 68.300 53.750 68.800 54.200 ;
        RECT 143.150 65.250 144.050 66.150 ;
        RECT 80.000 48.600 80.600 49.200 ;
        RECT 110.250 48.700 110.850 49.200 ;
        RECT 137.750 48.500 138.550 49.300 ;
        RECT 150.550 49.300 151.150 49.900 ;
        RECT 156.600 41.100 157.100 41.550 ;
        RECT 112.450 40.300 112.950 40.800 ;
        RECT 76.650 36.150 77.150 36.700 ;
        RECT 153.350 14.100 153.950 14.700 ;
        RECT 134.500 13.250 135.050 13.750 ;
      LAYER met3 ;
        RECT 109.155 114.250 140.650 145.250 ;
        RECT 68.250 53.725 68.850 54.225 ;
        RECT 79.900 48.500 80.700 95.150 ;
        RECT 109.155 82.050 140.650 113.050 ;
        RECT 85.550 81.425 86.100 81.925 ;
        RECT 81.850 78.725 82.350 79.425 ;
        RECT 81.855 52.950 106.350 76.950 ;
        RECT 109.155 49.850 140.650 80.850 ;
        RECT 143.100 65.225 144.100 66.175 ;
        RECT 110.200 48.675 110.900 49.225 ;
        RECT 137.700 48.475 138.600 49.325 ;
        RECT 150.500 49.275 151.200 49.925 ;
        RECT 112.400 40.275 113.000 40.825 ;
        RECT 76.600 36.700 77.200 36.725 ;
        RECT 76.600 36.100 90.900 36.700 ;
        RECT 90.300 34.200 90.900 36.100 ;
        RECT 122.155 15.700 153.650 46.700 ;
        RECT 156.550 41.075 157.150 41.575 ;
        RECT 153.300 14.075 154.000 14.725 ;
        RECT 134.450 13.225 135.100 13.775 ;
      LAYER via3 ;
        RECT 140.230 114.390 140.550 145.110 ;
        RECT 68.300 53.750 68.800 54.200 ;
        RECT 140.230 82.190 140.550 112.910 ;
        RECT 85.600 81.450 86.050 81.900 ;
        RECT 81.900 78.750 82.300 79.400 ;
        RECT 81.955 53.090 82.275 76.810 ;
        RECT 140.230 49.990 140.550 80.710 ;
        RECT 143.150 65.250 144.050 66.150 ;
        RECT 110.250 48.700 110.850 49.200 ;
        RECT 137.750 48.500 138.550 49.300 ;
        RECT 150.550 49.300 151.150 49.900 ;
        RECT 112.450 40.300 112.950 40.800 ;
        RECT 90.350 34.250 90.850 34.750 ;
        RECT 153.230 15.840 153.550 46.560 ;
        RECT 156.600 41.100 157.100 41.550 ;
        RECT 153.350 14.100 153.950 14.700 ;
        RECT 134.500 13.250 135.050 13.750 ;
      LAYER met4 ;
        RECT 124.395 144.555 124.915 145.500 ;
        RECT 139.995 145.190 140.515 145.500 ;
        RECT 109.850 114.945 139.460 144.555 ;
        RECT 124.395 112.355 124.915 114.945 ;
        RECT 139.995 114.310 140.630 145.190 ;
        RECT 139.995 112.990 140.515 114.310 ;
        RECT 109.850 82.745 139.460 112.355 ;
        RECT 81.850 76.890 82.350 79.450 ;
        RECT 81.850 76.750 82.355 76.890 ;
        RECT 68.240 1.000 68.840 54.260 ;
        RECT 81.875 53.010 82.355 76.750 ;
        RECT 85.550 76.255 86.100 81.950 ;
        RECT 124.395 80.155 124.915 82.745 ;
        RECT 139.995 82.110 140.630 112.990 ;
        RECT 139.995 80.790 140.515 82.110 ;
        RECT 83.045 53.645 105.655 76.255 ;
        RECT 109.850 50.545 139.460 80.155 ;
        RECT 139.995 66.200 140.630 80.790 ;
        RECT 139.995 65.200 144.100 66.200 ;
        RECT 110.150 48.600 110.950 50.545 ;
        RECT 124.395 49.600 124.915 50.545 ;
        RECT 137.650 48.400 138.650 50.545 ;
        RECT 139.995 49.910 140.630 65.200 ;
        RECT 139.995 49.600 140.515 49.910 ;
        RECT 150.450 46.005 151.250 50.000 ;
        RECT 90.325 1.000 90.915 34.825 ;
        RECT 112.400 1.000 113.000 40.850 ;
        RECT 122.850 16.395 152.460 46.005 ;
        RECT 153.150 16.000 153.630 46.640 ;
        RECT 156.550 41.630 157.150 41.650 ;
        RECT 156.550 41.050 157.160 41.630 ;
        RECT 153.150 15.700 153.650 16.000 ;
        RECT 153.150 15.200 153.850 15.700 ;
        RECT 153.350 14.705 153.850 15.200 ;
        RECT 153.345 14.095 153.955 14.705 ;
        RECT 134.450 11.900 135.100 13.800 ;
        RECT 134.480 1.000 135.080 11.900 ;
        RECT 156.560 3.575 157.160 41.050 ;
        RECT 156.570 1.000 157.155 3.575 ;
  END
END tt_um_edsonsilva17_ldo
END LIBRARY

