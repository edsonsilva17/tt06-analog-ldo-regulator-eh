** sch_path: /foss/designs/cobaia/xschem/diodo-I-V-pnp.sch
**.subckt diodo-I-V-pnp
XM1 GND GND net1 GND sky130_fd_pr__pfet_01v8_lvt L=0.35 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
VD D GND 0
.save i(vd)
VD1 D net1 0
.save i(vd1)
**** begin user architecture code

** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt




*.DC SRCname START STOP STEP

.control
save all
dc VD -1.8 1.8 0.01
plot i(vd1)
.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
