magic
tech sky130A
magscale 1 2
timestamp 1712843110
<< error_p >>
rect -70 3200 -10 9400
rect 10 3200 70 9400
rect -70 -3100 -10 3100
rect 10 -3100 70 3100
rect -70 -9400 -10 -3200
rect 10 -9400 70 -3200
<< metal3 >>
rect -6309 9372 -10 9400
rect -6309 3228 -94 9372
rect -30 3228 -10 9372
rect -6309 3200 -10 3228
rect 10 9372 6309 9400
rect 10 3228 6225 9372
rect 6289 3228 6309 9372
rect 10 3200 6309 3228
rect -6309 3072 -10 3100
rect -6309 -3072 -94 3072
rect -30 -3072 -10 3072
rect -6309 -3100 -10 -3072
rect 10 3072 6309 3100
rect 10 -3072 6225 3072
rect 6289 -3072 6309 3072
rect 10 -3100 6309 -3072
rect -6309 -3228 -10 -3200
rect -6309 -9372 -94 -3228
rect -30 -9372 -10 -3228
rect -6309 -9400 -10 -9372
rect 10 -3228 6309 -3200
rect 10 -9372 6225 -3228
rect 6289 -9372 6309 -3228
rect 10 -9400 6309 -9372
<< via3 >>
rect -94 3228 -30 9372
rect 6225 3228 6289 9372
rect -94 -3072 -30 3072
rect 6225 -3072 6289 3072
rect -94 -9372 -30 -3228
rect 6225 -9372 6289 -3228
<< mimcap >>
rect -6209 9260 -209 9300
rect -6209 3340 -6169 9260
rect -249 3340 -209 9260
rect -6209 3300 -209 3340
rect 110 9260 6110 9300
rect 110 3340 150 9260
rect 6070 3340 6110 9260
rect 110 3300 6110 3340
rect -6209 2960 -209 3000
rect -6209 -2960 -6169 2960
rect -249 -2960 -209 2960
rect -6209 -3000 -209 -2960
rect 110 2960 6110 3000
rect 110 -2960 150 2960
rect 6070 -2960 6110 2960
rect 110 -3000 6110 -2960
rect -6209 -3340 -209 -3300
rect -6209 -9260 -6169 -3340
rect -249 -9260 -209 -3340
rect -6209 -9300 -209 -9260
rect 110 -3340 6110 -3300
rect 110 -9260 150 -3340
rect 6070 -9260 6110 -3340
rect 110 -9300 6110 -9260
<< mimcapcontact >>
rect -6169 3340 -249 9260
rect 150 3340 6070 9260
rect -6169 -2960 -249 2960
rect 150 -2960 6070 2960
rect -6169 -9260 -249 -3340
rect 150 -9260 6070 -3340
<< metal4 >>
rect -3261 9261 -3157 9450
rect -141 9388 -37 9450
rect -141 9372 -14 9388
rect -6170 9260 -248 9261
rect -6170 3340 -6169 9260
rect -249 3340 -248 9260
rect -6170 3339 -248 3340
rect -3261 2961 -3157 3339
rect -141 3228 -94 9372
rect -30 3228 -14 9372
rect 3058 9261 3162 9450
rect 6178 9388 6282 9450
rect 6178 9372 6305 9388
rect 149 9260 6071 9261
rect 149 3340 150 9260
rect 6070 3340 6071 9260
rect 149 3339 6071 3340
rect -141 3212 -14 3228
rect -141 3088 -37 3212
rect -141 3072 -14 3088
rect -6170 2960 -248 2961
rect -6170 -2960 -6169 2960
rect -249 -2960 -248 2960
rect -6170 -2961 -248 -2960
rect -3261 -3339 -3157 -2961
rect -141 -3072 -94 3072
rect -30 -3072 -14 3072
rect 3058 2961 3162 3339
rect 6178 3228 6225 9372
rect 6289 3228 6305 9372
rect 6178 3212 6305 3228
rect 6178 3088 6282 3212
rect 6178 3072 6305 3088
rect 149 2960 6071 2961
rect 149 -2960 150 2960
rect 6070 -2960 6071 2960
rect 149 -2961 6071 -2960
rect -141 -3088 -14 -3072
rect -141 -3212 -37 -3088
rect -141 -3228 -14 -3212
rect -6170 -3340 -248 -3339
rect -6170 -9260 -6169 -3340
rect -249 -9260 -248 -3340
rect -6170 -9261 -248 -9260
rect -3261 -9450 -3157 -9261
rect -141 -9372 -94 -3228
rect -30 -9372 -14 -3228
rect 3058 -3339 3162 -2961
rect 6178 -3072 6225 3072
rect 6289 -3072 6305 3072
rect 6178 -3088 6305 -3072
rect 6178 -3212 6282 -3088
rect 6178 -3228 6305 -3212
rect 149 -3340 6071 -3339
rect 149 -9260 150 -3340
rect 6070 -9260 6071 -3340
rect 149 -9261 6071 -9260
rect -141 -9388 -14 -9372
rect -141 -9450 -37 -9388
rect 3058 -9450 3162 -9261
rect 6178 -9372 6225 -3228
rect 6289 -9372 6305 -3228
rect 6178 -9388 6305 -9372
rect 6178 -9450 6282 -9388
<< properties >>
string FIXED_BBOX 10 3200 6210 9400
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.0 l 30.0 val 1.822k carea 2.00 cperi 0.19 nx 2 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
