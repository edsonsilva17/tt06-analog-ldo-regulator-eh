magic
tech sky130A
magscale 1 2
timestamp 1713034554
<< metal1 >>
rect 0 10930 200 10950
rect 6020 10930 6220 10950
rect 0 10770 3240 10930
rect 0 10750 200 10770
rect 20 7860 180 10750
rect 3090 10290 3240 10770
rect 4660 10910 6220 10930
rect 4660 10790 5580 10910
rect 5700 10790 6220 10910
rect 4660 10770 6220 10790
rect 4660 10440 4810 10770
rect 6020 10750 6220 10770
rect 5000 10340 5720 10440
rect 3900 10120 4030 10200
rect 3900 10030 3920 10120
rect 4010 10030 4030 10120
rect 3900 10010 4030 10030
rect 20 7740 40 7860
rect 160 7740 180 7860
rect 20 7720 180 7740
rect 5560 4920 5720 10340
rect 5990 3600 6190 3620
rect 5740 3440 6190 3600
rect 5990 3420 6190 3440
rect 5790 3020 5950 3040
rect 5790 2910 5810 3020
rect 5930 2910 5950 3020
rect 30 2580 40 2700
rect 160 2580 170 2700
rect 5790 2590 5950 2910
rect 5990 2590 6190 2610
rect 5740 2430 6190 2590
rect 5990 2410 6190 2430
rect 5560 1730 5720 1750
rect 5560 1620 5580 1730
rect 5700 1620 5720 1730
rect 5560 1600 5720 1620
rect 20 700 180 950
rect 0 500 200 700
<< via1 >>
rect 5580 10790 5700 10910
rect 3920 10030 4010 10120
rect 40 7740 160 7860
rect 5810 2910 5930 3020
rect 40 2580 160 2700
rect 5580 1620 5700 1730
<< metal2 >>
rect 5580 10910 5700 10920
rect 5580 10780 5700 10790
rect 4030 10130 5950 10140
rect 3900 10120 5950 10130
rect 3900 10030 3920 10120
rect 4010 10030 5950 10120
rect 3900 10010 5950 10030
rect 20 7860 180 7880
rect 20 7740 40 7860
rect 160 7740 180 7860
rect 20 2700 180 7740
rect 5790 3020 5950 10010
rect 5790 2910 5810 3020
rect 5930 2910 5950 3020
rect 5790 2890 5950 2910
rect 20 2580 40 2700
rect 160 2580 180 2700
rect 20 2570 180 2580
rect 5580 1730 5700 1740
rect 5580 1610 5700 1620
<< via2 >>
rect 5580 10790 5700 10910
rect 5580 1620 5700 1730
<< metal3 >>
rect 5560 10910 5720 10930
rect 5560 10790 5580 10910
rect 5700 10790 5720 10910
rect 5560 1730 5720 10790
rect 5560 1620 5580 1730
rect 5700 1620 5720 1730
rect 5560 1600 5720 1620
use sky130_fd_pr__nfet_03v3_nvt_VP9Q5R  XM1
timestamp 1713034554
transform 0 1 3965 -1 0 10389
box -278 -1258 278 1258
use Ota_esq  x1
timestamp 1713034554
transform 1 0 170 0 1 4390
box -170 -3790 5570 5650
<< labels >>
flabel metal1 0 500 200 700 0 FreeSans 256 0 0 0 ldo_ibias
port 4 nsew
flabel metal1 0 10750 200 10950 0 FreeSans 256 0 0 0 ldo_in
port 1 nsew
flabel metal1 6020 10750 6220 10950 0 FreeSans 256 0 0 0 ldo_out
port 0 nsew
flabel metal1 5990 2410 6190 2610 0 FreeSans 256 0 0 0 ldo_gnd
port 2 nsew
flabel metal1 5990 3420 6190 3620 0 FreeSans 256 0 0 0 ldo_ref
port 3 nsew
<< end >>
