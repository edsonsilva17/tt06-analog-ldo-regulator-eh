magic
tech sky130A
magscale 1 2
timestamp 1712937985
<< pwell >>
rect -278 -1258 278 1258
<< nnmos >>
rect -50 -1000 50 1000
<< mvndiff >>
rect -108 988 -50 1000
rect -108 -988 -96 988
rect -62 -988 -50 988
rect -108 -1000 -50 -988
rect 50 988 108 1000
rect 50 -988 62 988
rect 96 -988 108 988
rect 50 -1000 108 -988
<< mvndiffc >>
rect -96 -988 -62 988
rect 62 -988 96 988
<< mvpsubdiff >>
rect -242 1210 242 1222
rect -242 1176 -134 1210
rect 134 1176 242 1210
rect -242 1164 242 1176
rect -242 1114 -184 1164
rect -242 -1114 -230 1114
rect -196 -1114 -184 1114
rect 184 1114 242 1164
rect -242 -1164 -184 -1114
rect 184 -1114 196 1114
rect 230 -1114 242 1114
rect 184 -1164 242 -1114
rect -242 -1176 242 -1164
rect -242 -1210 -134 -1176
rect 134 -1210 242 -1176
rect -242 -1222 242 -1210
<< mvpsubdiffcont >>
rect -134 1176 134 1210
rect -230 -1114 -196 1114
rect 196 -1114 230 1114
rect -134 -1210 134 -1176
<< poly >>
rect -50 1072 50 1088
rect -50 1038 -34 1072
rect 34 1038 50 1072
rect -50 1000 50 1038
rect -50 -1038 50 -1000
rect -50 -1072 -34 -1038
rect 34 -1072 50 -1038
rect -50 -1088 50 -1072
<< polycont >>
rect -34 1038 34 1072
rect -34 -1072 34 -1038
<< locali >>
rect -230 1176 -134 1210
rect 134 1176 230 1210
rect -230 1114 -196 1176
rect 196 1114 230 1176
rect -50 1038 -34 1072
rect 34 1038 50 1072
rect -96 988 -62 1004
rect -96 -1004 -62 -988
rect 62 988 96 1004
rect 62 -1004 96 -988
rect -50 -1072 -34 -1038
rect 34 -1072 50 -1038
rect -230 -1176 -196 -1114
rect 196 -1176 230 -1114
rect -230 -1210 -134 -1176
rect 134 -1210 230 -1176
<< viali >>
rect -34 1038 34 1072
rect -230 -176 -196 176
rect -96 -971 -62 -181
rect 62 181 96 971
rect -34 -1072 34 -1038
<< metal1 >>
rect -46 1072 46 1078
rect -46 1038 -34 1072
rect 34 1038 46 1072
rect -46 1032 46 1038
rect 56 971 102 983
rect -236 176 -190 188
rect -236 -176 -230 176
rect -196 -176 -190 176
rect 56 181 62 971
rect 96 181 102 971
rect 56 169 102 181
rect -236 -188 -190 -176
rect -102 -181 -56 -169
rect -102 -971 -96 -181
rect -62 -971 -56 -181
rect -102 -983 -56 -971
rect -46 -1038 46 -1032
rect -46 -1072 -34 -1038
rect 34 -1072 46 -1038
rect -46 -1078 46 -1072
<< properties >>
string FIXED_BBOX -213 -1193 213 1193
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 10.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -40 viadrn +40 viagate 100 viagb 0 viagr 0 viagl 15 viagt 0
<< end >>
