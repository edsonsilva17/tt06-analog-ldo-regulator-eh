magic
tech sky130A
magscale 1 2
timestamp 1712852575
<< nwell >>
rect -1906 -597 1906 597
<< mvpmos >>
rect -1648 -300 -1448 300
rect -1390 -300 -1190 300
rect -1132 -300 -932 300
rect -874 -300 -674 300
rect -616 -300 -416 300
rect -358 -300 -158 300
rect -100 -300 100 300
rect 158 -300 358 300
rect 416 -300 616 300
rect 674 -300 874 300
rect 932 -300 1132 300
rect 1190 -300 1390 300
rect 1448 -300 1648 300
<< mvpdiff >>
rect -1706 288 -1648 300
rect -1706 -288 -1694 288
rect -1660 -288 -1648 288
rect -1706 -300 -1648 -288
rect -1448 288 -1390 300
rect -1448 -288 -1436 288
rect -1402 -288 -1390 288
rect -1448 -300 -1390 -288
rect -1190 288 -1132 300
rect -1190 -288 -1178 288
rect -1144 -288 -1132 288
rect -1190 -300 -1132 -288
rect -932 288 -874 300
rect -932 -288 -920 288
rect -886 -288 -874 288
rect -932 -300 -874 -288
rect -674 288 -616 300
rect -674 -288 -662 288
rect -628 -288 -616 288
rect -674 -300 -616 -288
rect -416 288 -358 300
rect -416 -288 -404 288
rect -370 -288 -358 288
rect -416 -300 -358 -288
rect -158 288 -100 300
rect -158 -288 -146 288
rect -112 -288 -100 288
rect -158 -300 -100 -288
rect 100 288 158 300
rect 100 -288 112 288
rect 146 -288 158 288
rect 100 -300 158 -288
rect 358 288 416 300
rect 358 -288 370 288
rect 404 -288 416 288
rect 358 -300 416 -288
rect 616 288 674 300
rect 616 -288 628 288
rect 662 -288 674 288
rect 616 -300 674 -288
rect 874 288 932 300
rect 874 -288 886 288
rect 920 -288 932 288
rect 874 -300 932 -288
rect 1132 288 1190 300
rect 1132 -288 1144 288
rect 1178 -288 1190 288
rect 1132 -300 1190 -288
rect 1390 288 1448 300
rect 1390 -288 1402 288
rect 1436 -288 1448 288
rect 1390 -300 1448 -288
rect 1648 288 1706 300
rect 1648 -288 1660 288
rect 1694 -288 1706 288
rect 1648 -300 1706 -288
<< mvpdiffc >>
rect -1694 -288 -1660 288
rect -1436 -288 -1402 288
rect -1178 -288 -1144 288
rect -920 -288 -886 288
rect -662 -288 -628 288
rect -404 -288 -370 288
rect -146 -288 -112 288
rect 112 -288 146 288
rect 370 -288 404 288
rect 628 -288 662 288
rect 886 -288 920 288
rect 1144 -288 1178 288
rect 1402 -288 1436 288
rect 1660 -288 1694 288
<< mvnsubdiff >>
rect -1840 519 1840 531
rect -1840 485 -1732 519
rect 1732 485 1840 519
rect -1840 473 1840 485
rect -1840 423 -1782 473
rect -1840 -423 -1828 423
rect -1794 -423 -1782 423
rect 1782 423 1840 473
rect -1840 -473 -1782 -423
rect 1782 -423 1794 423
rect 1828 -423 1840 423
rect 1782 -473 1840 -423
rect -1840 -485 1840 -473
rect -1840 -519 -1732 -485
rect 1732 -519 1840 -485
rect -1840 -531 1840 -519
<< mvnsubdiffcont >>
rect -1732 485 1732 519
rect -1828 -423 -1794 423
rect 1794 -423 1828 423
rect -1732 -519 1732 -485
<< poly >>
rect -1648 381 -1448 397
rect -1648 347 -1632 381
rect -1464 347 -1448 381
rect -1648 300 -1448 347
rect -1390 381 -1190 397
rect -1390 347 -1374 381
rect -1206 347 -1190 381
rect -1390 300 -1190 347
rect -1132 381 -932 397
rect -1132 347 -1116 381
rect -948 347 -932 381
rect -1132 300 -932 347
rect -874 381 -674 397
rect -874 347 -858 381
rect -690 347 -674 381
rect -874 300 -674 347
rect -616 381 -416 397
rect -616 347 -600 381
rect -432 347 -416 381
rect -616 300 -416 347
rect -358 381 -158 397
rect -358 347 -342 381
rect -174 347 -158 381
rect -358 300 -158 347
rect -100 381 100 397
rect -100 347 -84 381
rect 84 347 100 381
rect -100 300 100 347
rect 158 381 358 397
rect 158 347 174 381
rect 342 347 358 381
rect 158 300 358 347
rect 416 381 616 397
rect 416 347 432 381
rect 600 347 616 381
rect 416 300 616 347
rect 674 381 874 397
rect 674 347 690 381
rect 858 347 874 381
rect 674 300 874 347
rect 932 381 1132 397
rect 932 347 948 381
rect 1116 347 1132 381
rect 932 300 1132 347
rect 1190 381 1390 397
rect 1190 347 1206 381
rect 1374 347 1390 381
rect 1190 300 1390 347
rect 1448 381 1648 397
rect 1448 347 1464 381
rect 1632 347 1648 381
rect 1448 300 1648 347
rect -1648 -347 -1448 -300
rect -1648 -381 -1632 -347
rect -1464 -381 -1448 -347
rect -1648 -397 -1448 -381
rect -1390 -347 -1190 -300
rect -1390 -381 -1374 -347
rect -1206 -381 -1190 -347
rect -1390 -397 -1190 -381
rect -1132 -347 -932 -300
rect -1132 -381 -1116 -347
rect -948 -381 -932 -347
rect -1132 -397 -932 -381
rect -874 -347 -674 -300
rect -874 -381 -858 -347
rect -690 -381 -674 -347
rect -874 -397 -674 -381
rect -616 -347 -416 -300
rect -616 -381 -600 -347
rect -432 -381 -416 -347
rect -616 -397 -416 -381
rect -358 -347 -158 -300
rect -358 -381 -342 -347
rect -174 -381 -158 -347
rect -358 -397 -158 -381
rect -100 -347 100 -300
rect -100 -381 -84 -347
rect 84 -381 100 -347
rect -100 -397 100 -381
rect 158 -347 358 -300
rect 158 -381 174 -347
rect 342 -381 358 -347
rect 158 -397 358 -381
rect 416 -347 616 -300
rect 416 -381 432 -347
rect 600 -381 616 -347
rect 416 -397 616 -381
rect 674 -347 874 -300
rect 674 -381 690 -347
rect 858 -381 874 -347
rect 674 -397 874 -381
rect 932 -347 1132 -300
rect 932 -381 948 -347
rect 1116 -381 1132 -347
rect 932 -397 1132 -381
rect 1190 -347 1390 -300
rect 1190 -381 1206 -347
rect 1374 -381 1390 -347
rect 1190 -397 1390 -381
rect 1448 -347 1648 -300
rect 1448 -381 1464 -347
rect 1632 -381 1648 -347
rect 1448 -397 1648 -381
<< polycont >>
rect -1632 347 -1464 381
rect -1374 347 -1206 381
rect -1116 347 -948 381
rect -858 347 -690 381
rect -600 347 -432 381
rect -342 347 -174 381
rect -84 347 84 381
rect 174 347 342 381
rect 432 347 600 381
rect 690 347 858 381
rect 948 347 1116 381
rect 1206 347 1374 381
rect 1464 347 1632 381
rect -1632 -381 -1464 -347
rect -1374 -381 -1206 -347
rect -1116 -381 -948 -347
rect -858 -381 -690 -347
rect -600 -381 -432 -347
rect -342 -381 -174 -347
rect -84 -381 84 -347
rect 174 -381 342 -347
rect 432 -381 600 -347
rect 690 -381 858 -347
rect 948 -381 1116 -347
rect 1206 -381 1374 -347
rect 1464 -381 1632 -347
<< locali >>
rect -1828 485 -1732 519
rect 1732 485 1828 519
rect 1794 423 1828 485
rect -1648 347 -1632 381
rect -1464 347 -1448 381
rect -1390 347 -1374 381
rect -1206 347 -1190 381
rect -1132 347 -1116 381
rect -948 347 -932 381
rect -874 347 -858 381
rect -690 347 -674 381
rect -616 347 -600 381
rect -432 347 -416 381
rect -358 347 -342 381
rect -174 347 -158 381
rect -100 347 -84 381
rect 84 347 100 381
rect 158 347 174 381
rect 342 347 358 381
rect 416 347 432 381
rect 600 347 616 381
rect 674 347 690 381
rect 858 347 874 381
rect 932 347 948 381
rect 1116 347 1132 381
rect 1190 347 1206 381
rect 1374 347 1390 381
rect 1448 347 1464 381
rect 1632 347 1648 381
rect -1694 288 -1660 304
rect -1694 -304 -1660 -288
rect -1436 288 -1402 304
rect -1436 -304 -1402 -288
rect -1178 288 -1144 304
rect -1178 -304 -1144 -288
rect -920 288 -886 304
rect -920 -304 -886 -288
rect -662 288 -628 304
rect -662 -304 -628 -288
rect -404 288 -370 304
rect -404 -304 -370 -288
rect -146 288 -112 304
rect -146 -304 -112 -288
rect 112 288 146 304
rect 112 -304 146 -288
rect 370 288 404 304
rect 370 -304 404 -288
rect 628 288 662 304
rect 628 -304 662 -288
rect 886 288 920 304
rect 886 -304 920 -288
rect 1144 288 1178 304
rect 1144 -304 1178 -288
rect 1402 288 1436 304
rect 1402 -304 1436 -288
rect 1660 288 1694 304
rect 1660 -304 1694 -288
rect -1648 -381 -1632 -347
rect -1464 -381 -1448 -347
rect -1390 -381 -1374 -347
rect -1206 -381 -1190 -347
rect -1132 -381 -1116 -347
rect -948 -381 -932 -347
rect -874 -381 -858 -347
rect -690 -381 -674 -347
rect -616 -381 -600 -347
rect -432 -381 -416 -347
rect -358 -381 -342 -347
rect -174 -381 -158 -347
rect -100 -381 -84 -347
rect 84 -381 100 -347
rect 158 -381 174 -347
rect 342 -381 358 -347
rect 416 -381 432 -347
rect 600 -381 616 -347
rect 674 -381 690 -347
rect 858 -381 874 -347
rect 932 -381 948 -347
rect 1116 -381 1132 -347
rect 1190 -381 1206 -347
rect 1374 -381 1390 -347
rect 1448 -381 1464 -347
rect 1632 -381 1648 -347
rect -1828 -485 -1794 -423
rect 1794 -485 1828 -423
rect -1828 -519 -1732 -485
rect 1732 -519 1828 -485
<< viali >>
rect -1828 423 -1794 485
rect -1828 97 -1794 423
rect -1632 347 -1464 381
rect -1374 347 -1206 381
rect -1116 347 -948 381
rect -858 347 -690 381
rect -600 347 -432 381
rect -342 347 -174 381
rect -84 347 84 381
rect 174 347 342 381
rect 432 347 600 381
rect 690 347 858 381
rect 948 347 1116 381
rect 1206 347 1374 381
rect 1464 347 1632 381
rect -1694 41 -1660 271
rect -1436 -271 -1402 -41
rect -1178 41 -1144 271
rect -920 -271 -886 -41
rect -662 41 -628 271
rect -404 -271 -370 -41
rect -146 41 -112 271
rect 112 -271 146 -41
rect 370 41 404 271
rect 628 -271 662 -41
rect 886 41 920 271
rect 1144 -271 1178 -41
rect 1402 41 1436 271
rect 1660 -271 1694 -41
rect -1632 -381 -1464 -347
rect -1374 -381 -1206 -347
rect -1116 -381 -948 -347
rect -858 -381 -690 -347
rect -600 -381 -432 -347
rect -342 -381 -174 -347
rect -84 -381 84 -347
rect 174 -381 342 -347
rect 432 -381 600 -347
rect 690 -381 858 -347
rect 948 -381 1116 -347
rect 1206 -381 1374 -347
rect 1464 -381 1632 -347
<< metal1 >>
rect -1834 485 -1788 497
rect -1834 97 -1828 485
rect -1794 97 -1788 485
rect -1644 381 -1452 387
rect -1644 347 -1632 381
rect -1464 347 -1452 381
rect -1644 341 -1452 347
rect -1386 381 -1194 387
rect -1386 347 -1374 381
rect -1206 347 -1194 381
rect -1386 341 -1194 347
rect -1128 381 -936 387
rect -1128 347 -1116 381
rect -948 347 -936 381
rect -1128 341 -936 347
rect -870 381 -678 387
rect -870 347 -858 381
rect -690 347 -678 381
rect -870 341 -678 347
rect -612 381 -420 387
rect -612 347 -600 381
rect -432 347 -420 381
rect -612 341 -420 347
rect -354 381 -162 387
rect -354 347 -342 381
rect -174 347 -162 381
rect -354 341 -162 347
rect -96 381 96 387
rect -96 347 -84 381
rect 84 347 96 381
rect -96 341 96 347
rect 162 381 354 387
rect 162 347 174 381
rect 342 347 354 381
rect 162 341 354 347
rect 420 381 612 387
rect 420 347 432 381
rect 600 347 612 381
rect 420 341 612 347
rect 678 381 870 387
rect 678 347 690 381
rect 858 347 870 381
rect 678 341 870 347
rect 936 381 1128 387
rect 936 347 948 381
rect 1116 347 1128 381
rect 936 341 1128 347
rect 1194 381 1386 387
rect 1194 347 1206 381
rect 1374 347 1386 381
rect 1194 341 1386 347
rect 1452 381 1644 387
rect 1452 347 1464 381
rect 1632 347 1644 381
rect 1452 341 1644 347
rect -1834 85 -1788 97
rect -1700 271 -1654 283
rect -1700 41 -1694 271
rect -1660 41 -1654 271
rect -1700 29 -1654 41
rect -1184 271 -1138 283
rect -1184 41 -1178 271
rect -1144 41 -1138 271
rect -1184 29 -1138 41
rect -668 271 -622 283
rect -668 41 -662 271
rect -628 41 -622 271
rect -668 29 -622 41
rect -152 271 -106 283
rect -152 41 -146 271
rect -112 41 -106 271
rect -152 29 -106 41
rect 364 271 410 283
rect 364 41 370 271
rect 404 41 410 271
rect 364 29 410 41
rect 880 271 926 283
rect 880 41 886 271
rect 920 41 926 271
rect 880 29 926 41
rect 1396 271 1442 283
rect 1396 41 1402 271
rect 1436 41 1442 271
rect 1396 29 1442 41
rect -1442 -41 -1396 -29
rect -1442 -271 -1436 -41
rect -1402 -271 -1396 -41
rect -1442 -283 -1396 -271
rect -926 -41 -880 -29
rect -926 -271 -920 -41
rect -886 -271 -880 -41
rect -926 -283 -880 -271
rect -410 -41 -364 -29
rect -410 -271 -404 -41
rect -370 -271 -364 -41
rect -410 -283 -364 -271
rect 106 -41 152 -29
rect 106 -271 112 -41
rect 146 -271 152 -41
rect 106 -283 152 -271
rect 622 -41 668 -29
rect 622 -271 628 -41
rect 662 -271 668 -41
rect 622 -283 668 -271
rect 1138 -41 1184 -29
rect 1138 -271 1144 -41
rect 1178 -271 1184 -41
rect 1138 -283 1184 -271
rect 1654 -41 1700 -29
rect 1654 -271 1660 -41
rect 1694 -271 1700 -41
rect 1654 -283 1700 -271
rect -1644 -347 -1452 -341
rect -1644 -381 -1632 -347
rect -1464 -381 -1452 -347
rect -1644 -387 -1452 -381
rect -1386 -347 -1194 -341
rect -1386 -381 -1374 -347
rect -1206 -381 -1194 -347
rect -1386 -387 -1194 -381
rect -1128 -347 -936 -341
rect -1128 -381 -1116 -347
rect -948 -381 -936 -347
rect -1128 -387 -936 -381
rect -870 -347 -678 -341
rect -870 -381 -858 -347
rect -690 -381 -678 -347
rect -870 -387 -678 -381
rect -612 -347 -420 -341
rect -612 -381 -600 -347
rect -432 -381 -420 -347
rect -612 -387 -420 -381
rect -354 -347 -162 -341
rect -354 -381 -342 -347
rect -174 -381 -162 -347
rect -354 -387 -162 -381
rect -96 -347 96 -341
rect -96 -381 -84 -347
rect 84 -381 96 -347
rect -96 -387 96 -381
rect 162 -347 354 -341
rect 162 -381 174 -347
rect 342 -381 354 -347
rect 162 -387 354 -381
rect 420 -347 612 -341
rect 420 -381 432 -347
rect 600 -381 612 -347
rect 420 -387 612 -381
rect 678 -347 870 -341
rect 678 -381 690 -347
rect 858 -381 870 -347
rect 678 -387 870 -381
rect 936 -347 1128 -341
rect 936 -381 948 -347
rect 1116 -381 1128 -347
rect 936 -387 1128 -381
rect 1194 -347 1386 -341
rect 1194 -381 1206 -347
rect 1374 -381 1386 -347
rect 1194 -387 1386 -381
rect 1452 -347 1644 -341
rect 1452 -381 1464 -347
rect 1632 -381 1644 -347
rect 1452 -387 1644 -381
<< properties >>
string FIXED_BBOX -1811 -502 1811 502
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 3.0 l 1.0 m 1 nf 13 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl -40 viagt 0
<< end >>
