magic
tech sky130A
magscale 1 2
timestamp 1712795588
<< metal3 >>
rect -3150 34572 3149 34600
rect -3150 28428 3065 34572
rect 3129 28428 3149 34572
rect -3150 28400 3149 28428
rect -3150 28272 3149 28300
rect -3150 22128 3065 28272
rect 3129 22128 3149 28272
rect -3150 22100 3149 22128
rect -3150 21972 3149 22000
rect -3150 15828 3065 21972
rect 3129 15828 3149 21972
rect -3150 15800 3149 15828
rect -3150 15672 3149 15700
rect -3150 9528 3065 15672
rect 3129 9528 3149 15672
rect -3150 9500 3149 9528
rect -3150 9372 3149 9400
rect -3150 3228 3065 9372
rect 3129 3228 3149 9372
rect -3150 3200 3149 3228
rect -3150 3072 3149 3100
rect -3150 -3072 3065 3072
rect 3129 -3072 3149 3072
rect -3150 -3100 3149 -3072
rect -3150 -3228 3149 -3200
rect -3150 -9372 3065 -3228
rect 3129 -9372 3149 -3228
rect -3150 -9400 3149 -9372
rect -3150 -9528 3149 -9500
rect -3150 -15672 3065 -9528
rect 3129 -15672 3149 -9528
rect -3150 -15700 3149 -15672
rect -3150 -15828 3149 -15800
rect -3150 -21972 3065 -15828
rect 3129 -21972 3149 -15828
rect -3150 -22000 3149 -21972
rect -3150 -22128 3149 -22100
rect -3150 -28272 3065 -22128
rect 3129 -28272 3149 -22128
rect -3150 -28300 3149 -28272
rect -3150 -28428 3149 -28400
rect -3150 -34572 3065 -28428
rect 3129 -34572 3149 -28428
rect -3150 -34600 3149 -34572
<< via3 >>
rect 3065 28428 3129 34572
rect 3065 22128 3129 28272
rect 3065 15828 3129 21972
rect 3065 9528 3129 15672
rect 3065 3228 3129 9372
rect 3065 -3072 3129 3072
rect 3065 -9372 3129 -3228
rect 3065 -15672 3129 -9528
rect 3065 -21972 3129 -15828
rect 3065 -28272 3129 -22128
rect 3065 -34572 3129 -28428
<< mimcap >>
rect -3050 34460 2950 34500
rect -3050 28540 -3010 34460
rect 2910 28540 2950 34460
rect -3050 28500 2950 28540
rect -3050 28160 2950 28200
rect -3050 22240 -3010 28160
rect 2910 22240 2950 28160
rect -3050 22200 2950 22240
rect -3050 21860 2950 21900
rect -3050 15940 -3010 21860
rect 2910 15940 2950 21860
rect -3050 15900 2950 15940
rect -3050 15560 2950 15600
rect -3050 9640 -3010 15560
rect 2910 9640 2950 15560
rect -3050 9600 2950 9640
rect -3050 9260 2950 9300
rect -3050 3340 -3010 9260
rect 2910 3340 2950 9260
rect -3050 3300 2950 3340
rect -3050 2960 2950 3000
rect -3050 -2960 -3010 2960
rect 2910 -2960 2950 2960
rect -3050 -3000 2950 -2960
rect -3050 -3340 2950 -3300
rect -3050 -9260 -3010 -3340
rect 2910 -9260 2950 -3340
rect -3050 -9300 2950 -9260
rect -3050 -9640 2950 -9600
rect -3050 -15560 -3010 -9640
rect 2910 -15560 2950 -9640
rect -3050 -15600 2950 -15560
rect -3050 -15940 2950 -15900
rect -3050 -21860 -3010 -15940
rect 2910 -21860 2950 -15940
rect -3050 -21900 2950 -21860
rect -3050 -22240 2950 -22200
rect -3050 -28160 -3010 -22240
rect 2910 -28160 2950 -22240
rect -3050 -28200 2950 -28160
rect -3050 -28540 2950 -28500
rect -3050 -34460 -3010 -28540
rect 2910 -34460 2950 -28540
rect -3050 -34500 2950 -34460
<< mimcapcontact >>
rect -3010 28540 2910 34460
rect -3010 22240 2910 28160
rect -3010 15940 2910 21860
rect -3010 9640 2910 15560
rect -3010 3340 2910 9260
rect -3010 -2960 2910 2960
rect -3010 -9260 2910 -3340
rect -3010 -15560 2910 -9640
rect -3010 -21860 2910 -15940
rect -3010 -28160 2910 -22240
rect -3010 -34460 2910 -28540
<< metal4 >>
rect -102 34461 2 34650
rect 3018 34588 3122 34650
rect 3018 34572 3145 34588
rect -3011 34460 2911 34461
rect -3011 28540 -3010 34460
rect 2910 28540 2911 34460
rect -3011 28539 2911 28540
rect -102 28161 2 28539
rect 3018 28428 3065 34572
rect 3129 28428 3145 34572
rect 3018 28412 3145 28428
rect 3018 28288 3122 28412
rect 3018 28272 3145 28288
rect -3011 28160 2911 28161
rect -3011 22240 -3010 28160
rect 2910 22240 2911 28160
rect -3011 22239 2911 22240
rect -102 21861 2 22239
rect 3018 22128 3065 28272
rect 3129 22128 3145 28272
rect 3018 22112 3145 22128
rect 3018 21988 3122 22112
rect 3018 21972 3145 21988
rect -3011 21860 2911 21861
rect -3011 15940 -3010 21860
rect 2910 15940 2911 21860
rect -3011 15939 2911 15940
rect -102 15561 2 15939
rect 3018 15828 3065 21972
rect 3129 15828 3145 21972
rect 3018 15812 3145 15828
rect 3018 15688 3122 15812
rect 3018 15672 3145 15688
rect -3011 15560 2911 15561
rect -3011 9640 -3010 15560
rect 2910 9640 2911 15560
rect -3011 9639 2911 9640
rect -102 9261 2 9639
rect 3018 9528 3065 15672
rect 3129 9528 3145 15672
rect 3018 9512 3145 9528
rect 3018 9388 3122 9512
rect 3018 9372 3145 9388
rect -3011 9260 2911 9261
rect -3011 3340 -3010 9260
rect 2910 3340 2911 9260
rect -3011 3339 2911 3340
rect -102 2961 2 3339
rect 3018 3228 3065 9372
rect 3129 3228 3145 9372
rect 3018 3212 3145 3228
rect 3018 3088 3122 3212
rect 3018 3072 3145 3088
rect -3011 2960 2911 2961
rect -3011 -2960 -3010 2960
rect 2910 -2960 2911 2960
rect -3011 -2961 2911 -2960
rect -102 -3339 2 -2961
rect 3018 -3072 3065 3072
rect 3129 -3072 3145 3072
rect 3018 -3088 3145 -3072
rect 3018 -3212 3122 -3088
rect 3018 -3228 3145 -3212
rect -3011 -3340 2911 -3339
rect -3011 -9260 -3010 -3340
rect 2910 -9260 2911 -3340
rect -3011 -9261 2911 -9260
rect -102 -9639 2 -9261
rect 3018 -9372 3065 -3228
rect 3129 -9372 3145 -3228
rect 3018 -9388 3145 -9372
rect 3018 -9512 3122 -9388
rect 3018 -9528 3145 -9512
rect -3011 -9640 2911 -9639
rect -3011 -15560 -3010 -9640
rect 2910 -15560 2911 -9640
rect -3011 -15561 2911 -15560
rect -102 -15939 2 -15561
rect 3018 -15672 3065 -9528
rect 3129 -15672 3145 -9528
rect 3018 -15688 3145 -15672
rect 3018 -15812 3122 -15688
rect 3018 -15828 3145 -15812
rect -3011 -15940 2911 -15939
rect -3011 -21860 -3010 -15940
rect 2910 -21860 2911 -15940
rect -3011 -21861 2911 -21860
rect -102 -22239 2 -21861
rect 3018 -21972 3065 -15828
rect 3129 -21972 3145 -15828
rect 3018 -21988 3145 -21972
rect 3018 -22112 3122 -21988
rect 3018 -22128 3145 -22112
rect -3011 -22240 2911 -22239
rect -3011 -28160 -3010 -22240
rect 2910 -28160 2911 -22240
rect -3011 -28161 2911 -28160
rect -102 -28539 2 -28161
rect 3018 -28272 3065 -22128
rect 3129 -28272 3145 -22128
rect 3018 -28288 3145 -28272
rect 3018 -28412 3122 -28288
rect 3018 -28428 3145 -28412
rect -3011 -28540 2911 -28539
rect -3011 -34460 -3010 -28540
rect 2910 -34460 2911 -28540
rect -3011 -34461 2911 -34460
rect -102 -34650 2 -34461
rect 3018 -34572 3065 -28428
rect 3129 -34572 3145 -28428
rect 3018 -34588 3145 -34572
rect 3018 -34650 3122 -34588
<< properties >>
string FIXED_BBOX -3150 28400 3050 34600
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.0 l 30.0 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 11 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
