magic
tech sky130A
magscale 1 2
timestamp 1712930560
<< pwell >>
rect -1102 -558 1102 558
<< mvnmos >>
rect -874 -300 -674 300
rect -616 -300 -416 300
rect -358 -300 -158 300
rect -100 -300 100 300
rect 158 -300 358 300
rect 416 -300 616 300
rect 674 -300 874 300
<< mvndiff >>
rect -932 288 -874 300
rect -932 -288 -920 288
rect -886 -288 -874 288
rect -932 -300 -874 -288
rect -674 288 -616 300
rect -674 -288 -662 288
rect -628 -288 -616 288
rect -674 -300 -616 -288
rect -416 288 -358 300
rect -416 -288 -404 288
rect -370 -288 -358 288
rect -416 -300 -358 -288
rect -158 288 -100 300
rect -158 -288 -146 288
rect -112 -288 -100 288
rect -158 -300 -100 -288
rect 100 288 158 300
rect 100 -288 112 288
rect 146 -288 158 288
rect 100 -300 158 -288
rect 358 288 416 300
rect 358 -288 370 288
rect 404 -288 416 288
rect 358 -300 416 -288
rect 616 288 674 300
rect 616 -288 628 288
rect 662 -288 674 288
rect 616 -300 674 -288
rect 874 288 932 300
rect 874 -288 886 288
rect 920 -288 932 288
rect 874 -300 932 -288
<< mvndiffc >>
rect -920 -288 -886 288
rect -662 -288 -628 288
rect -404 -288 -370 288
rect -146 -288 -112 288
rect 112 -288 146 288
rect 370 -288 404 288
rect 628 -288 662 288
rect 886 -288 920 288
<< mvpsubdiff >>
rect -1066 510 1066 522
rect -1066 476 -958 510
rect 958 476 1066 510
rect -1066 464 1066 476
rect -1066 414 -1008 464
rect -1066 -414 -1054 414
rect -1020 -414 -1008 414
rect 1008 414 1066 464
rect -1066 -464 -1008 -414
rect 1008 -414 1020 414
rect 1054 -414 1066 414
rect 1008 -464 1066 -414
rect -1066 -476 1066 -464
rect -1066 -510 -958 -476
rect 958 -510 1066 -476
rect -1066 -522 1066 -510
<< mvpsubdiffcont >>
rect -958 476 958 510
rect -1054 -414 -1020 414
rect 1020 -414 1054 414
rect -958 -510 958 -476
<< poly >>
rect -874 372 -674 388
rect -874 338 -858 372
rect -690 338 -674 372
rect -874 300 -674 338
rect -616 372 -416 388
rect -616 338 -600 372
rect -432 338 -416 372
rect -616 300 -416 338
rect -358 372 -158 388
rect -358 338 -342 372
rect -174 338 -158 372
rect -358 300 -158 338
rect -100 372 100 388
rect -100 338 -84 372
rect 84 338 100 372
rect -100 300 100 338
rect 158 372 358 388
rect 158 338 174 372
rect 342 338 358 372
rect 158 300 358 338
rect 416 372 616 388
rect 416 338 432 372
rect 600 338 616 372
rect 416 300 616 338
rect 674 372 874 388
rect 674 338 690 372
rect 858 338 874 372
rect 674 300 874 338
rect -874 -338 -674 -300
rect -874 -372 -858 -338
rect -690 -372 -674 -338
rect -874 -388 -674 -372
rect -616 -338 -416 -300
rect -616 -372 -600 -338
rect -432 -372 -416 -338
rect -616 -388 -416 -372
rect -358 -338 -158 -300
rect -358 -372 -342 -338
rect -174 -372 -158 -338
rect -358 -388 -158 -372
rect -100 -338 100 -300
rect -100 -372 -84 -338
rect 84 -372 100 -338
rect -100 -388 100 -372
rect 158 -338 358 -300
rect 158 -372 174 -338
rect 342 -372 358 -338
rect 158 -388 358 -372
rect 416 -338 616 -300
rect 416 -372 432 -338
rect 600 -372 616 -338
rect 416 -388 616 -372
rect 674 -338 874 -300
rect 674 -372 690 -338
rect 858 -372 874 -338
rect 674 -388 874 -372
<< polycont >>
rect -858 338 -690 372
rect -600 338 -432 372
rect -342 338 -174 372
rect -84 338 84 372
rect 174 338 342 372
rect 432 338 600 372
rect 690 338 858 372
rect -858 -372 -690 -338
rect -600 -372 -432 -338
rect -342 -372 -174 -338
rect -84 -372 84 -338
rect 174 -372 342 -338
rect 432 -372 600 -338
rect 690 -372 858 -338
<< locali >>
rect -1054 476 -958 510
rect 958 476 1054 510
rect -1054 414 -1020 476
rect 1020 414 1054 476
rect -874 338 -858 372
rect -690 338 -674 372
rect -616 338 -600 372
rect -432 338 -416 372
rect -358 338 -342 372
rect -174 338 -158 372
rect -100 338 -84 372
rect 84 338 100 372
rect 158 338 174 372
rect 342 338 358 372
rect 416 338 432 372
rect 600 338 616 372
rect 674 338 690 372
rect 858 338 874 372
rect -920 288 -886 304
rect -920 -304 -886 -288
rect -662 288 -628 304
rect -662 -304 -628 -288
rect -404 288 -370 304
rect -404 -304 -370 -288
rect -146 288 -112 304
rect -146 -304 -112 -288
rect 112 288 146 304
rect 112 -304 146 -288
rect 370 288 404 304
rect 370 -304 404 -288
rect 628 288 662 304
rect 628 -304 662 -288
rect 886 288 920 304
rect 886 -304 920 -288
rect -874 -372 -858 -338
rect -690 -372 -674 -338
rect -616 -372 -600 -338
rect -432 -372 -416 -338
rect -358 -372 -342 -338
rect -174 -372 -158 -338
rect -100 -372 -84 -338
rect 84 -372 100 -338
rect 158 -372 174 -338
rect 342 -372 358 -338
rect 416 -372 432 -338
rect 600 -372 616 -338
rect 674 -372 690 -338
rect 858 -372 874 -338
rect 1020 -476 1054 -414
rect -1054 -510 -958 -476
rect 958 -510 1054 -476
<< viali >>
rect -858 338 -690 372
rect -600 338 -432 372
rect -342 338 -174 372
rect -84 338 84 372
rect 174 338 342 372
rect 432 338 600 372
rect 690 338 858 372
rect -1054 -414 -1020 0
rect -920 41 -886 271
rect -662 -271 -628 -41
rect -404 41 -370 271
rect -146 -271 -112 -41
rect 112 41 146 271
rect 370 -271 404 -41
rect 628 41 662 271
rect 886 -271 920 -41
rect -858 -372 -690 -338
rect -600 -372 -432 -338
rect -342 -372 -174 -338
rect -84 -372 84 -338
rect 174 -372 342 -338
rect 432 -372 600 -338
rect 690 -372 858 -338
rect -1054 -476 -1020 -414
<< metal1 >>
rect -870 372 -678 378
rect -870 338 -858 372
rect -690 338 -678 372
rect -870 332 -678 338
rect -612 372 -420 378
rect -612 338 -600 372
rect -432 338 -420 372
rect -612 332 -420 338
rect -354 372 -162 378
rect -354 338 -342 372
rect -174 338 -162 372
rect -354 332 -162 338
rect -96 372 96 378
rect -96 338 -84 372
rect 84 338 96 372
rect -96 332 96 338
rect 162 372 354 378
rect 162 338 174 372
rect 342 338 354 372
rect 162 332 354 338
rect 420 372 612 378
rect 420 338 432 372
rect 600 338 612 372
rect 420 332 612 338
rect 678 372 870 378
rect 678 338 690 372
rect 858 338 870 372
rect 678 332 870 338
rect -926 271 -880 283
rect -926 41 -920 271
rect -886 41 -880 271
rect -926 29 -880 41
rect -410 271 -364 283
rect -410 41 -404 271
rect -370 41 -364 271
rect -410 29 -364 41
rect 106 271 152 283
rect 106 41 112 271
rect 146 41 152 271
rect 106 29 152 41
rect 622 271 668 283
rect 622 41 628 271
rect 662 41 668 271
rect 622 29 668 41
rect -1060 0 -1014 12
rect -1060 -476 -1054 0
rect -1020 -476 -1014 0
rect -668 -41 -622 -29
rect -668 -271 -662 -41
rect -628 -271 -622 -41
rect -668 -283 -622 -271
rect -152 -41 -106 -29
rect -152 -271 -146 -41
rect -112 -271 -106 -41
rect -152 -283 -106 -271
rect 364 -41 410 -29
rect 364 -271 370 -41
rect 404 -271 410 -41
rect 364 -283 410 -271
rect 880 -41 926 -29
rect 880 -271 886 -41
rect 920 -271 926 -41
rect 880 -283 926 -271
rect -870 -338 -678 -332
rect -870 -372 -858 -338
rect -690 -372 -678 -338
rect -870 -378 -678 -372
rect -612 -338 -420 -332
rect -612 -372 -600 -338
rect -432 -372 -420 -338
rect -612 -378 -420 -372
rect -354 -338 -162 -332
rect -354 -372 -342 -338
rect -174 -372 -162 -338
rect -354 -378 -162 -372
rect -96 -338 96 -332
rect -96 -372 -84 -338
rect 84 -372 96 -338
rect -96 -378 96 -372
rect 162 -338 354 -332
rect 162 -372 174 -338
rect 342 -372 354 -338
rect 162 -378 354 -372
rect 420 -338 612 -332
rect 420 -372 432 -338
rect 600 -372 612 -338
rect 420 -378 612 -372
rect 678 -338 870 -332
rect 678 -372 690 -338
rect 858 -372 870 -338
rect 678 -378 870 -372
rect -1060 -488 -1014 -476
<< properties >>
string FIXED_BBOX -1037 -493 1037 493
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3.0 l 1.0 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl +50 viagt 0
<< end >>
