magic
tech sky130A
magscale 1 2
timestamp 1713034554
<< metal1 >>
rect 5370 500 5570 530
rect -150 490 5570 500
rect -150 360 5070 490
rect 5150 360 5570 490
rect -150 350 5570 360
rect -150 -710 10 350
rect 5370 330 5570 350
rect 1580 170 5550 190
rect 1580 60 5410 170
rect 5530 60 5550 170
rect 1580 40 5550 60
rect 4310 -60 4320 -50
rect 1770 -130 4320 -60
rect 4310 -140 4320 -130
rect 4410 -140 4420 -50
rect -150 -860 3280 -710
rect 5370 -820 5570 -770
rect 4410 -920 5570 -820
rect -150 -1180 3540 -1030
rect 4410 -1180 4510 -920
rect 5370 -970 5570 -920
rect -150 -1310 40 -1180
rect -150 -2110 10 -1310
rect 190 -1360 3490 -1270
rect 1040 -1650 1130 -1360
rect 3980 -1500 4390 -1350
rect 4520 -1370 5040 -1350
rect 4520 -1480 4750 -1370
rect 4860 -1480 5040 -1370
rect 4520 -1500 5040 -1480
rect 5160 -1370 5550 -1350
rect 5160 -1480 5410 -1370
rect 5530 -1480 5550 -1370
rect 5160 -1500 5550 -1480
rect 1040 -1660 3490 -1650
rect 1040 -1730 1050 -1660
rect 1120 -1730 3490 -1660
rect 1040 -1740 3490 -1730
rect 3980 -1830 4210 -1500
rect 1430 -1980 4210 -1830
rect 5050 -1850 5150 -1660
rect 5390 -1780 5550 -1500
rect -170 -2140 30 -2110
rect -170 -2290 3274 -2140
rect 3980 -2270 4210 -1980
rect 4750 -1910 5150 -1850
rect 4750 -2270 4850 -1910
rect 5050 -2100 5150 -1910
rect 5370 -1980 5570 -1780
rect 5390 -2270 5550 -1980
rect -170 -2310 30 -2290
rect -150 -2960 10 -2310
rect 3980 -2420 4390 -2270
rect 4520 -2420 5040 -2270
rect 5160 -2420 5550 -2270
rect 4410 -2840 4510 -2580
rect 5370 -2840 5570 -2790
rect 4410 -2940 5570 -2840
rect -150 -3110 3534 -2960
rect 5370 -2990 5570 -2940
rect -170 -3270 30 -3240
rect -170 -3300 3280 -3270
rect -170 -3390 1040 -3300
rect 1130 -3390 3280 -3300
rect -170 -3420 3280 -3390
rect -170 -3440 30 -3420
rect 1040 -3510 1130 -3420
rect 1040 -3600 3490 -3510
<< via1 >>
rect 5070 360 5150 490
rect 5410 60 5530 170
rect 4320 -140 4410 -50
rect 4750 -1480 4860 -1370
rect 5410 -1480 5530 -1370
rect 1050 -1730 1120 -1660
rect 1040 -3390 1130 -3300
<< metal2 >>
rect 5070 490 5150 500
rect 5070 350 5150 360
rect 5390 170 5550 190
rect 5390 60 5410 170
rect 5530 60 5550 170
rect 4310 -50 4420 -40
rect 4310 -140 4320 -50
rect 4410 -140 4420 -50
rect 4310 -660 4420 -140
rect 4310 -770 4860 -660
rect 4750 -1370 4860 -770
rect 4750 -1490 4860 -1480
rect 5390 -1370 5550 60
rect 5390 -1480 5410 -1370
rect 5530 -1480 5550 -1370
rect 5390 -1500 5550 -1480
rect 1040 -1660 1130 -1650
rect 1040 -1730 1050 -1660
rect 1120 -1730 1130 -1660
rect 1040 -3300 1130 -1730
rect 1040 -3400 1130 -3390
<< via2 >>
rect 5070 360 5150 490
rect 4320 -140 4410 -50
<< metal3 >>
rect 5060 490 5160 495
rect 5060 360 5070 490
rect 5150 360 5160 490
rect 5060 355 5160 360
rect 4310 -50 4420 -45
rect 4310 -140 4320 -50
rect 4410 -140 4420 -50
rect 4310 -145 4420 -140
<< via3 >>
rect 5070 360 5150 490
rect 4320 -140 4410 -50
<< metal4 >>
rect 4310 -50 4420 1110
rect 5060 490 5160 890
rect 5060 360 5070 490
rect 5150 360 5160 490
rect 5060 350 5160 360
rect 4310 -140 4320 -50
rect 4410 -140 4420 -50
rect 4310 -150 4420 -140
use sky130_fd_pr__cap_mim_m3_1_M5BWMD  XC1
timestamp 1713034554
transform 1 0 2710 0 1 3250
box -2450 -2400 2449 2400
use sky130_fd_pr__pfet_g5v0d10v5_4LQ75H  XM1
timestamp 1713034554
transform -1 0 4458 0 -1 -2343
box -308 -497 308 497
use sky130_fd_pr__pfet_g5v0d10v5_LMT75H  XM2
timestamp 1713034554
transform 1 0 4458 0 1 -1423
box -308 -497 308 497
use sky130_fd_pr__nfet_g5v0d10v5_RVNTYK  XM3
timestamp 1713034554
transform -1 0 5100 0 -1 -2830
box -278 -958 278 958
use sky130_fd_pr__nfet_g5v0d10v5_RMPAXK  XM4
timestamp 1713034554
transform 1 0 5100 0 1 -930
box -278 -958 278 958
use sky130_fd_pr__pfet_g5v0d10v5_FYUU4F  XM5
timestamp 1713034554
transform 1 0 2481 0 1 -2063
box -1261 -597 1261 597
use sky130_fd_pr__pfet_g5v0d10v5_C5553C  XM6
timestamp 1713034554
transform 1 0 1836 0 1 -943
box -1906 -597 1906 597
use sky130_fd_pr__nfet_g5v0d10v5_YCT7Q3  XM7
timestamp 1713034554
transform 1 0 2644 0 1 270
box -1102 -558 1102 558
use sky130_fd_pr__pfet_g5v0d10v5_FY4V4F  XM8
timestamp 1713034554
transform 1 0 2481 0 1 -3193
box -1261 -597 1261 597
<< labels >>
flabel metal1 -170 -2310 30 -2110 0 FreeSans 256 0 0 0 VDD
port 2 nsew
flabel metal1 -170 -3440 30 -3240 0 FreeSans 256 0 0 0 Ibias
port 4 nsew
flabel metal1 5370 -1980 5570 -1780 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 5370 330 5570 530 0 FreeSans 256 0 0 0 Vout
port 5 nsew
flabel metal1 5370 -970 5570 -770 0 FreeSans 256 0 0 0 Vip
port 1 nsew
flabel metal1 5370 -2990 5570 -2790 0 FreeSans 256 0 0 0 Vin
port 0 nsew
<< end >>
