magic
tech sky130A
magscale 1 2
timestamp 1712944184
<< error_p >>
rect -287 881 -225 887
rect -159 881 -97 887
rect -31 881 31 887
rect 97 881 159 887
rect 225 881 287 887
rect -287 847 -275 881
rect -159 847 -147 881
rect -31 847 -19 881
rect 97 847 109 881
rect 225 847 237 881
rect -287 841 -225 847
rect -159 841 -97 847
rect -31 841 31 847
rect 97 841 159 847
rect 225 841 287 847
rect -287 -847 -225 -841
rect -159 -847 -97 -841
rect -31 -847 31 -841
rect 97 -847 159 -841
rect 225 -847 287 -841
rect -287 -881 -275 -847
rect -159 -881 -147 -847
rect -31 -881 -19 -847
rect 97 -881 109 -847
rect 225 -881 237 -847
rect -287 -887 -225 -881
rect -159 -887 -97 -881
rect -31 -887 31 -881
rect 97 -887 159 -881
rect 225 -887 287 -881
<< nwell >>
rect -487 -1019 487 1019
<< pmoslvt >>
rect -291 -800 -221 800
rect -163 -800 -93 800
rect -35 -800 35 800
rect 93 -800 163 800
rect 221 -800 291 800
<< pdiff >>
rect -349 788 -291 800
rect -349 -788 -337 788
rect -303 -788 -291 788
rect -349 -800 -291 -788
rect -221 788 -163 800
rect -221 -788 -209 788
rect -175 -788 -163 788
rect -221 -800 -163 -788
rect -93 788 -35 800
rect -93 -788 -81 788
rect -47 -788 -35 788
rect -93 -800 -35 -788
rect 35 788 93 800
rect 35 -788 47 788
rect 81 -788 93 788
rect 35 -800 93 -788
rect 163 788 221 800
rect 163 -788 175 788
rect 209 -788 221 788
rect 163 -800 221 -788
rect 291 788 349 800
rect 291 -788 303 788
rect 337 -788 349 788
rect 291 -800 349 -788
<< pdiffc >>
rect -337 -788 -303 788
rect -209 -788 -175 788
rect -81 -788 -47 788
rect 47 -788 81 788
rect 175 -788 209 788
rect 303 -788 337 788
<< nsubdiff >>
rect -451 949 -355 983
rect 355 949 451 983
rect -451 887 -417 949
rect 417 887 451 949
rect -451 -949 -417 -887
rect 417 -949 451 -887
rect -451 -983 -355 -949
rect 355 -983 451 -949
<< nsubdiffcont >>
rect -355 949 355 983
rect -451 -887 -417 887
rect 417 -887 451 887
rect -355 -983 355 -949
<< poly >>
rect -291 881 -221 897
rect -291 847 -275 881
rect -237 847 -221 881
rect -291 800 -221 847
rect -163 881 -93 897
rect -163 847 -147 881
rect -109 847 -93 881
rect -163 800 -93 847
rect -35 881 35 897
rect -35 847 -19 881
rect 19 847 35 881
rect -35 800 35 847
rect 93 881 163 897
rect 93 847 109 881
rect 147 847 163 881
rect 93 800 163 847
rect 221 881 291 897
rect 221 847 237 881
rect 275 847 291 881
rect 221 800 291 847
rect -291 -847 -221 -800
rect -291 -881 -275 -847
rect -237 -881 -221 -847
rect -291 -897 -221 -881
rect -163 -847 -93 -800
rect -163 -881 -147 -847
rect -109 -881 -93 -847
rect -163 -897 -93 -881
rect -35 -847 35 -800
rect -35 -881 -19 -847
rect 19 -881 35 -847
rect -35 -897 35 -881
rect 93 -847 163 -800
rect 93 -881 109 -847
rect 147 -881 163 -847
rect 93 -897 163 -881
rect 221 -847 291 -800
rect 221 -881 237 -847
rect 275 -881 291 -847
rect 221 -897 291 -881
<< polycont >>
rect -275 847 -237 881
rect -147 847 -109 881
rect -19 847 19 881
rect 109 847 147 881
rect 237 847 275 881
rect -275 -881 -237 -847
rect -147 -881 -109 -847
rect -19 -881 19 -847
rect 109 -881 147 -847
rect 237 -881 275 -847
<< locali >>
rect -451 949 -355 983
rect 355 949 451 983
rect -451 887 -417 949
rect 417 887 451 949
rect -291 847 -275 881
rect -237 847 -221 881
rect -163 847 -147 881
rect -109 847 -93 881
rect -35 847 -19 881
rect 19 847 35 881
rect 93 847 109 881
rect 147 847 163 881
rect 221 847 237 881
rect 275 847 291 881
rect -337 788 -303 804
rect -337 -804 -303 -788
rect -209 788 -175 804
rect -209 -804 -175 -788
rect -81 788 -47 804
rect -81 -804 -47 -788
rect 47 788 81 804
rect 47 -804 81 -788
rect 175 788 209 804
rect 175 -804 209 -788
rect 303 788 337 804
rect 303 -804 337 -788
rect -291 -881 -275 -847
rect -237 -881 -221 -847
rect -163 -881 -147 -847
rect -109 -881 -93 -847
rect -35 -881 -19 -847
rect 19 -881 35 -847
rect 93 -881 109 -847
rect 147 -881 163 -847
rect 221 -881 237 -847
rect 275 -881 291 -847
rect -451 -949 -417 -887
rect 417 -949 451 -887
rect -451 -983 -355 -949
rect 355 -983 451 -949
<< viali >>
rect -208 949 208 983
rect -275 847 -237 881
rect -147 847 -109 881
rect -19 847 19 881
rect 109 847 147 881
rect 237 847 275 881
rect -337 141 -303 771
rect -209 -771 -175 -141
rect -81 141 -47 771
rect 47 -771 81 -141
rect 175 141 209 771
rect 303 -771 337 -141
rect -275 -881 -237 -847
rect -147 -881 -109 -847
rect -19 -881 19 -847
rect 109 -881 147 -847
rect 237 -881 275 -847
<< metal1 >>
rect -220 983 220 989
rect -220 949 -208 983
rect 208 949 220 983
rect -220 943 220 949
rect -287 881 -225 887
rect -287 847 -275 881
rect -237 847 -225 881
rect -287 841 -225 847
rect -159 881 -97 887
rect -159 847 -147 881
rect -109 847 -97 881
rect -159 841 -97 847
rect -31 881 31 887
rect -31 847 -19 881
rect 19 847 31 881
rect -31 841 31 847
rect 97 881 159 887
rect 97 847 109 881
rect 147 847 159 881
rect 97 841 159 847
rect 225 881 287 887
rect 225 847 237 881
rect 275 847 287 881
rect 225 841 287 847
rect -343 771 -297 783
rect -343 141 -337 771
rect -303 141 -297 771
rect -343 129 -297 141
rect -87 771 -41 783
rect -87 141 -81 771
rect -47 141 -41 771
rect -87 129 -41 141
rect 169 771 215 783
rect 169 141 175 771
rect 209 141 215 771
rect 169 129 215 141
rect -215 -141 -169 -129
rect -215 -771 -209 -141
rect -175 -771 -169 -141
rect -215 -783 -169 -771
rect 41 -141 87 -129
rect 41 -771 47 -141
rect 81 -771 87 -141
rect 41 -783 87 -771
rect 297 -141 343 -129
rect 297 -771 303 -141
rect 337 -771 343 -141
rect 297 -783 343 -771
rect -287 -847 -225 -841
rect -287 -881 -275 -847
rect -237 -881 -225 -847
rect -287 -887 -225 -881
rect -159 -847 -97 -841
rect -159 -881 -147 -847
rect -109 -881 -97 -847
rect -159 -887 -97 -881
rect -31 -847 31 -841
rect -31 -881 -19 -847
rect 19 -881 31 -847
rect -31 -887 31 -881
rect 97 -847 159 -841
rect 97 -881 109 -847
rect 147 -881 159 -847
rect 97 -887 159 -881
rect 225 -847 287 -841
rect 225 -881 237 -847
rect 275 -881 287 -847
rect 225 -887 287 -881
<< properties >>
string FIXED_BBOX -434 -966 434 966
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 8.0 l 0.35 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 50
<< end >>
