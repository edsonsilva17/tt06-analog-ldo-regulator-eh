magic
tech sky130A
magscale 1 2
timestamp 1712843110
<< error_p >>
rect -3230 6350 -3170 12550
rect -3150 6350 -3090 12550
rect 3089 6350 3149 12550
rect 3169 6350 3229 12550
rect -3230 50 -3170 6250
rect -3150 50 -3090 6250
rect 3089 50 3149 6250
rect 3169 50 3229 6250
rect -3230 -6250 -3170 -50
rect -3150 -6250 -3090 -50
rect 3089 -6250 3149 -50
rect 3169 -6250 3229 -50
rect -3230 -12550 -3170 -6350
rect -3150 -12550 -3090 -6350
rect 3089 -12550 3149 -6350
rect 3169 -12550 3229 -6350
<< metal3 >>
rect -9469 12522 -3170 12550
rect -9469 6378 -3254 12522
rect -3190 6378 -3170 12522
rect -9469 6350 -3170 6378
rect -3150 12522 3149 12550
rect -3150 6378 3065 12522
rect 3129 6378 3149 12522
rect -3150 6350 3149 6378
rect 3169 12522 9468 12550
rect 3169 6378 9384 12522
rect 9448 6378 9468 12522
rect 3169 6350 9468 6378
rect -9469 6222 -3170 6250
rect -9469 78 -3254 6222
rect -3190 78 -3170 6222
rect -9469 50 -3170 78
rect -3150 6222 3149 6250
rect -3150 78 3065 6222
rect 3129 78 3149 6222
rect -3150 50 3149 78
rect 3169 6222 9468 6250
rect 3169 78 9384 6222
rect 9448 78 9468 6222
rect 3169 50 9468 78
rect -9469 -78 -3170 -50
rect -9469 -6222 -3254 -78
rect -3190 -6222 -3170 -78
rect -9469 -6250 -3170 -6222
rect -3150 -78 3149 -50
rect -3150 -6222 3065 -78
rect 3129 -6222 3149 -78
rect -3150 -6250 3149 -6222
rect 3169 -78 9468 -50
rect 3169 -6222 9384 -78
rect 9448 -6222 9468 -78
rect 3169 -6250 9468 -6222
rect -9469 -6378 -3170 -6350
rect -9469 -12522 -3254 -6378
rect -3190 -12522 -3170 -6378
rect -9469 -12550 -3170 -12522
rect -3150 -6378 3149 -6350
rect -3150 -12522 3065 -6378
rect 3129 -12522 3149 -6378
rect -3150 -12550 3149 -12522
rect 3169 -6378 9468 -6350
rect 3169 -12522 9384 -6378
rect 9448 -12522 9468 -6378
rect 3169 -12550 9468 -12522
<< via3 >>
rect -3254 6378 -3190 12522
rect 3065 6378 3129 12522
rect 9384 6378 9448 12522
rect -3254 78 -3190 6222
rect 3065 78 3129 6222
rect 9384 78 9448 6222
rect -3254 -6222 -3190 -78
rect 3065 -6222 3129 -78
rect 9384 -6222 9448 -78
rect -3254 -12522 -3190 -6378
rect 3065 -12522 3129 -6378
rect 9384 -12522 9448 -6378
<< mimcap >>
rect -9369 12410 -3369 12450
rect -9369 6490 -9329 12410
rect -3409 6490 -3369 12410
rect -9369 6450 -3369 6490
rect -3050 12410 2950 12450
rect -3050 6490 -3010 12410
rect 2910 6490 2950 12410
rect -3050 6450 2950 6490
rect 3269 12410 9269 12450
rect 3269 6490 3309 12410
rect 9229 6490 9269 12410
rect 3269 6450 9269 6490
rect -9369 6110 -3369 6150
rect -9369 190 -9329 6110
rect -3409 190 -3369 6110
rect -9369 150 -3369 190
rect -3050 6110 2950 6150
rect -3050 190 -3010 6110
rect 2910 190 2950 6110
rect -3050 150 2950 190
rect 3269 6110 9269 6150
rect 3269 190 3309 6110
rect 9229 190 9269 6110
rect 3269 150 9269 190
rect -9369 -190 -3369 -150
rect -9369 -6110 -9329 -190
rect -3409 -6110 -3369 -190
rect -9369 -6150 -3369 -6110
rect -3050 -190 2950 -150
rect -3050 -6110 -3010 -190
rect 2910 -6110 2950 -190
rect -3050 -6150 2950 -6110
rect 3269 -190 9269 -150
rect 3269 -6110 3309 -190
rect 9229 -6110 9269 -190
rect 3269 -6150 9269 -6110
rect -9369 -6490 -3369 -6450
rect -9369 -12410 -9329 -6490
rect -3409 -12410 -3369 -6490
rect -9369 -12450 -3369 -12410
rect -3050 -6490 2950 -6450
rect -3050 -12410 -3010 -6490
rect 2910 -12410 2950 -6490
rect -3050 -12450 2950 -12410
rect 3269 -6490 9269 -6450
rect 3269 -12410 3309 -6490
rect 9229 -12410 9269 -6490
rect 3269 -12450 9269 -12410
<< mimcapcontact >>
rect -9329 6490 -3409 12410
rect -3010 6490 2910 12410
rect 3309 6490 9229 12410
rect -9329 190 -3409 6110
rect -3010 190 2910 6110
rect 3309 190 9229 6110
rect -9329 -6110 -3409 -190
rect -3010 -6110 2910 -190
rect 3309 -6110 9229 -190
rect -9329 -12410 -3409 -6490
rect -3010 -12410 2910 -6490
rect 3309 -12410 9229 -6490
<< metal4 >>
rect -6421 12411 -6317 12600
rect -3301 12538 -3197 12600
rect -3301 12522 -3174 12538
rect -9330 12410 -3408 12411
rect -9330 6490 -9329 12410
rect -3409 6490 -3408 12410
rect -9330 6489 -3408 6490
rect -6421 6111 -6317 6489
rect -3301 6378 -3254 12522
rect -3190 6378 -3174 12522
rect -102 12411 2 12600
rect 3018 12538 3122 12600
rect 3018 12522 3145 12538
rect -3011 12410 2911 12411
rect -3011 6490 -3010 12410
rect 2910 6490 2911 12410
rect -3011 6489 2911 6490
rect -3301 6362 -3174 6378
rect -3301 6238 -3197 6362
rect -3301 6222 -3174 6238
rect -9330 6110 -3408 6111
rect -9330 190 -9329 6110
rect -3409 190 -3408 6110
rect -9330 189 -3408 190
rect -6421 -189 -6317 189
rect -3301 78 -3254 6222
rect -3190 78 -3174 6222
rect -102 6111 2 6489
rect 3018 6378 3065 12522
rect 3129 6378 3145 12522
rect 6217 12411 6321 12600
rect 9337 12538 9441 12600
rect 9337 12522 9464 12538
rect 3308 12410 9230 12411
rect 3308 6490 3309 12410
rect 9229 6490 9230 12410
rect 3308 6489 9230 6490
rect 3018 6362 3145 6378
rect 3018 6238 3122 6362
rect 3018 6222 3145 6238
rect -3011 6110 2911 6111
rect -3011 190 -3010 6110
rect 2910 190 2911 6110
rect -3011 189 2911 190
rect -3301 62 -3174 78
rect -3301 -62 -3197 62
rect -3301 -78 -3174 -62
rect -9330 -190 -3408 -189
rect -9330 -6110 -9329 -190
rect -3409 -6110 -3408 -190
rect -9330 -6111 -3408 -6110
rect -6421 -6489 -6317 -6111
rect -3301 -6222 -3254 -78
rect -3190 -6222 -3174 -78
rect -102 -189 2 189
rect 3018 78 3065 6222
rect 3129 78 3145 6222
rect 6217 6111 6321 6489
rect 9337 6378 9384 12522
rect 9448 6378 9464 12522
rect 9337 6362 9464 6378
rect 9337 6238 9441 6362
rect 9337 6222 9464 6238
rect 3308 6110 9230 6111
rect 3308 190 3309 6110
rect 9229 190 9230 6110
rect 3308 189 9230 190
rect 3018 62 3145 78
rect 3018 -62 3122 62
rect 3018 -78 3145 -62
rect -3011 -190 2911 -189
rect -3011 -6110 -3010 -190
rect 2910 -6110 2911 -190
rect -3011 -6111 2911 -6110
rect -3301 -6238 -3174 -6222
rect -3301 -6362 -3197 -6238
rect -3301 -6378 -3174 -6362
rect -9330 -6490 -3408 -6489
rect -9330 -12410 -9329 -6490
rect -3409 -12410 -3408 -6490
rect -9330 -12411 -3408 -12410
rect -6421 -12600 -6317 -12411
rect -3301 -12522 -3254 -6378
rect -3190 -12522 -3174 -6378
rect -102 -6489 2 -6111
rect 3018 -6222 3065 -78
rect 3129 -6222 3145 -78
rect 6217 -189 6321 189
rect 9337 78 9384 6222
rect 9448 78 9464 6222
rect 9337 62 9464 78
rect 9337 -62 9441 62
rect 9337 -78 9464 -62
rect 3308 -190 9230 -189
rect 3308 -6110 3309 -190
rect 9229 -6110 9230 -190
rect 3308 -6111 9230 -6110
rect 3018 -6238 3145 -6222
rect 3018 -6362 3122 -6238
rect 3018 -6378 3145 -6362
rect -3011 -6490 2911 -6489
rect -3011 -12410 -3010 -6490
rect 2910 -12410 2911 -6490
rect -3011 -12411 2911 -12410
rect -3301 -12538 -3174 -12522
rect -3301 -12600 -3197 -12538
rect -102 -12600 2 -12411
rect 3018 -12522 3065 -6378
rect 3129 -12522 3145 -6378
rect 6217 -6489 6321 -6111
rect 9337 -6222 9384 -78
rect 9448 -6222 9464 -78
rect 9337 -6238 9464 -6222
rect 9337 -6362 9441 -6238
rect 9337 -6378 9464 -6362
rect 3308 -6490 9230 -6489
rect 3308 -12410 3309 -6490
rect 9229 -12410 9230 -6490
rect 3308 -12411 9230 -12410
rect 3018 -12538 3145 -12522
rect 3018 -12600 3122 -12538
rect 6217 -12600 6321 -12411
rect 9337 -12522 9384 -6378
rect 9448 -12522 9464 -6378
rect 9337 -12538 9464 -12522
rect 9337 -12600 9441 -12538
<< properties >>
string FIXED_BBOX 3169 6350 9369 12550
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.0 l 30.0 val 1.822k carea 2.00 cperi 0.19 nx 3 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
