magic
tech sky130A
magscale 1 2
timestamp 1713034554
<< metal3 >>
rect -3150 9372 3149 9400
rect -3150 3228 3065 9372
rect 3129 3228 3149 9372
rect -3150 3200 3149 3228
rect -3150 2932 3149 2960
rect -3150 -3212 3065 2932
rect 3129 -3212 3149 2932
rect -3150 -3240 3149 -3212
rect -3150 -3508 3149 -3480
rect -3150 -9652 3065 -3508
rect 3129 -9652 3149 -3508
rect -3150 -9680 3149 -9652
<< via3 >>
rect 3065 3228 3129 9372
rect 3065 -3212 3129 2932
rect 3065 -9652 3129 -3508
<< mimcap >>
rect -3050 9260 2950 9300
rect -3050 3340 -3010 9260
rect 2910 3340 2950 9260
rect -3050 3300 2950 3340
rect -3050 2820 2950 2860
rect -3050 -3100 -3010 2820
rect 2910 -3100 2950 2820
rect -3050 -3140 2950 -3100
rect -3050 -3620 2950 -3580
rect -3050 -9540 -3010 -3620
rect 2910 -9540 2950 -3620
rect -3050 -9580 2950 -9540
<< mimcapcontact >>
rect -3010 3340 2910 9260
rect -3010 -3100 2910 2820
rect -3010 -9540 2910 -3620
<< metal4 >>
rect -102 9261 2 9450
rect 3018 9388 3122 9450
rect 3018 9372 3145 9388
rect -3011 9260 2911 9261
rect -3011 3340 -3010 9260
rect 2910 3340 2911 9260
rect -3011 3339 2911 3340
rect -102 2821 2 3339
rect 3018 3228 3065 9372
rect 3129 3228 3145 9372
rect 3018 3212 3145 3228
rect 3018 2948 3122 3212
rect 3018 2932 3145 2948
rect -3011 2820 2911 2821
rect -3011 -3100 -3010 2820
rect 2910 -3100 2911 2820
rect -3011 -3101 2911 -3100
rect -102 -3619 2 -3101
rect 3018 -3212 3065 2932
rect 3129 -3212 3145 2932
rect 3018 -3228 3145 -3212
rect 3018 -3492 3122 -3228
rect 3018 -3508 3145 -3492
rect -3011 -3620 2911 -3619
rect -3011 -9540 -3010 -3620
rect 2910 -9540 2911 -3620
rect -3011 -9541 2911 -9540
rect -102 -9730 2 -9541
rect 3018 -9652 3065 -3508
rect 3129 -9652 3145 -3508
rect 3018 -9668 3145 -9652
rect 3018 -9730 3122 -9668
<< properties >>
string FIXED_BBOX -3150 3200 3050 9400
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.0 l 30.0 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
